
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-32.95,39.6893,61.95,-63.2229</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>14.5,-13</position>
<gparam>LABEL_TEXT Go to https://cedar.to/vjyQw7 to download the latest version!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>14.5,-9.5</position>
<gparam>LABEL_TEXT Error: This file was made with a newer version of Cedar Logic!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 0>
</circuit>
<throw_away></throw_away>

	<version>2.3.5 | 2018-09-25 23:06:05</version><circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-191.804,22.75,177.129,-163.375</PageViewport>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>34.5,14</position>
<input>
<ID>IN_0</ID>491 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>0,-17.5</position>
<gparam>LABEL_TEXT Address Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>38.5,-118</position>
<input>
<ID>IN_0</ID>587 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID inc_tr</lparam></gate>
<gate>
<ID>2</ID>
<type>AI_RAM_12x16</type>
<position>23,12.5</position>
<input>
<ID>ADDRESS_0</ID>197 </input>
<input>
<ID>ADDRESS_1</ID>198 </input>
<input>
<ID>ADDRESS_10</ID>203 </input>
<input>
<ID>ADDRESS_11</ID>204 </input>
<input>
<ID>ADDRESS_2</ID>195 </input>
<input>
<ID>ADDRESS_3</ID>201 </input>
<input>
<ID>ADDRESS_4</ID>199 </input>
<input>
<ID>ADDRESS_5</ID>202 </input>
<input>
<ID>ADDRESS_6</ID>200 </input>
<input>
<ID>ADDRESS_7</ID>193 </input>
<input>
<ID>ADDRESS_8</ID>194 </input>
<input>
<ID>ADDRESS_9</ID>196 </input>
<input>
<ID>DATA_IN_0</ID>6 </input>
<input>
<ID>DATA_IN_1</ID>7 </input>
<input>
<ID>DATA_IN_10</ID>13 </input>
<input>
<ID>DATA_IN_11</ID>15 </input>
<input>
<ID>DATA_IN_12</ID>10 </input>
<input>
<ID>DATA_IN_13</ID>9 </input>
<input>
<ID>DATA_IN_14</ID>12 </input>
<input>
<ID>DATA_IN_15</ID>17 </input>
<input>
<ID>DATA_IN_2</ID>2 </input>
<input>
<ID>DATA_IN_3</ID>3 </input>
<input>
<ID>DATA_IN_4</ID>4 </input>
<input>
<ID>DATA_IN_5</ID>8 </input>
<input>
<ID>DATA_IN_6</ID>5 </input>
<input>
<ID>DATA_IN_7</ID>11 </input>
<input>
<ID>DATA_IN_8</ID>16 </input>
<input>
<ID>DATA_IN_9</ID>14 </input>
<output>
<ID>DATA_OUT_0</ID>6 </output>
<output>
<ID>DATA_OUT_1</ID>7 </output>
<output>
<ID>DATA_OUT_10</ID>13 </output>
<output>
<ID>DATA_OUT_11</ID>15 </output>
<output>
<ID>DATA_OUT_12</ID>10 </output>
<output>
<ID>DATA_OUT_13</ID>9 </output>
<output>
<ID>DATA_OUT_14</ID>12 </output>
<output>
<ID>DATA_OUT_15</ID>17 </output>
<output>
<ID>DATA_OUT_2</ID>2 </output>
<output>
<ID>DATA_OUT_3</ID>3 </output>
<output>
<ID>DATA_OUT_4</ID>4 </output>
<output>
<ID>DATA_OUT_5</ID>8 </output>
<output>
<ID>DATA_OUT_6</ID>5 </output>
<output>
<ID>DATA_OUT_7</ID>11 </output>
<output>
<ID>DATA_OUT_8</ID>16 </output>
<output>
<ID>DATA_OUT_9</ID>14 </output>
<input>
<ID>ENABLE_0</ID>564 </input>
<input>
<ID>write_clock</ID>491 </input>
<input>
<ID>write_enable</ID>563 </input>
<gparam>angle 0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam></gate>
<gate>
<ID>76</ID>
<type>DE_TO</type>
<position>-7,4.5</position>
<input>
<ID>IN_0</ID>492 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>12</ID>
<type>AI_REGISTER12</type>
<position>40,-53</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>107 </input>
<input>
<ID>IN_10</ID>106 </input>
<input>
<ID>IN_11</ID>101 </input>
<input>
<ID>IN_2</ID>109 </input>
<input>
<ID>IN_3</ID>110 </input>
<input>
<ID>IN_4</ID>99 </input>
<input>
<ID>IN_5</ID>104 </input>
<input>
<ID>IN_6</ID>105 </input>
<input>
<ID>IN_7</ID>100 </input>
<input>
<ID>IN_8</ID>103 </input>
<input>
<ID>IN_9</ID>102 </input>
<output>
<ID>OUT_0</ID>552 </output>
<output>
<ID>OUT_1</ID>557 </output>
<output>
<ID>OUT_10</ID>561 </output>
<output>
<ID>OUT_11</ID>562 </output>
<output>
<ID>OUT_2</ID>551 </output>
<output>
<ID>OUT_3</ID>556 </output>
<output>
<ID>OUT_4</ID>553 </output>
<output>
<ID>OUT_5</ID>554 </output>
<output>
<ID>OUT_6</ID>555 </output>
<output>
<ID>OUT_7</ID>558 </output>
<output>
<ID>OUT_8</ID>559 </output>
<output>
<ID>OUT_9</ID>560 </output>
<input>
<ID>clear</ID>569 </input>
<input>
<ID>clock</ID>498 </input>
<input>
<ID>count_enable</ID>572 </input>
<input>
<ID>count_up</ID>571 </input>
<input>
<ID>load</ID>570 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>39.5,-144.5</position>
<input>
<ID>IN_0</ID>589 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clr_tr</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_REGISTER8</type>
<position>3.5,-148.5</position>
<input>
<ID>IN_0</ID>609 </input>
<input>
<ID>IN_1</ID>610 </input>
<input>
<ID>IN_2</ID>611 </input>
<input>
<ID>IN_3</ID>614 </input>
<input>
<ID>IN_4</ID>615 </input>
<input>
<ID>IN_5</ID>616 </input>
<input>
<ID>IN_6</ID>612 </input>
<input>
<ID>IN_7</ID>613 </input>
<input>
<ID>clock</ID>493 </input>
<input>
<ID>count_up</ID>581 </input>
<input>
<ID>load</ID>591 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>0,-141</position>
<input>
<ID>IN_0</ID>591 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_or</lparam></gate>
<gate>
<ID>6</ID>
<type>AI_REGISTER12</type>
<position>-1,-31.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>179 </input>
<input>
<ID>IN_10</ID>177 </input>
<input>
<ID>IN_11</ID>178 </input>
<input>
<ID>IN_2</ID>93 </input>
<input>
<ID>IN_3</ID>96 </input>
<input>
<ID>IN_4</ID>97 </input>
<input>
<ID>IN_5</ID>98 </input>
<input>
<ID>IN_6</ID>176 </input>
<input>
<ID>IN_7</ID>94 </input>
<input>
<ID>IN_8</ID>180 </input>
<input>
<ID>IN_9</ID>175 </input>
<output>
<ID>OUT_0</ID>188 </output>
<output>
<ID>OUT_1</ID>182 </output>
<output>
<ID>OUT_10</ID>191 </output>
<output>
<ID>OUT_11</ID>192 </output>
<output>
<ID>OUT_2</ID>190 </output>
<output>
<ID>OUT_3</ID>189 </output>
<output>
<ID>OUT_4</ID>181 </output>
<output>
<ID>OUT_5</ID>183 </output>
<output>
<ID>OUT_6</ID>184 </output>
<output>
<ID>OUT_7</ID>185 </output>
<output>
<ID>OUT_8</ID>187 </output>
<output>
<ID>OUT_9</ID>186 </output>
<input>
<ID>clear</ID>565 </input>
<input>
<ID>clock</ID>499 </input>
<input>
<ID>count_enable</ID>568 </input>
<input>
<ID>load</ID>566 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>14</ID>
<type>AM_REGISTER16</type>
<position>36,-90</position>
<input>
<ID>IN_0</ID>254 </input>
<input>
<ID>IN_1</ID>255 </input>
<input>
<ID>IN_10</ID>261 </input>
<input>
<ID>IN_11</ID>266 </input>
<input>
<ID>IN_12</ID>262 </input>
<input>
<ID>IN_13</ID>265 </input>
<input>
<ID>IN_14</ID>263 </input>
<input>
<ID>IN_15</ID>264 </input>
<input>
<ID>IN_2</ID>256 </input>
<input>
<ID>IN_3</ID>257 </input>
<input>
<ID>IN_4</ID>258 </input>
<input>
<ID>IN_5</ID>269 </input>
<input>
<ID>IN_6</ID>259 </input>
<input>
<ID>IN_7</ID>268 </input>
<input>
<ID>IN_8</ID>260 </input>
<input>
<ID>IN_9</ID>267 </input>
<output>
<ID>OUT_0</ID>414 </output>
<output>
<ID>OUT_1</ID>399 </output>
<output>
<ID>OUT_10</ID>405 </output>
<output>
<ID>OUT_11</ID>403 </output>
<output>
<ID>OUT_12</ID>404 </output>
<output>
<ID>OUT_13</ID>406 </output>
<output>
<ID>OUT_14</ID>407 </output>
<output>
<ID>OUT_15</ID>409 </output>
<output>
<ID>OUT_2</ID>410 </output>
<output>
<ID>OUT_3</ID>400 </output>
<output>
<ID>OUT_4</ID>401 </output>
<output>
<ID>OUT_5</ID>408 </output>
<output>
<ID>OUT_6</ID>411 </output>
<output>
<ID>OUT_7</ID>412 </output>
<output>
<ID>OUT_8</ID>402 </output>
<output>
<ID>OUT_9</ID>413 </output>
<input>
<ID>clear</ID>583 </input>
<input>
<ID>clock</ID>496 </input>
<input>
<ID>count_enable</ID>577 </input>
<input>
<ID>count_up</ID>578 </input>
<input>
<ID>load</ID>582 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>-1,-158</position>
<input>
<ID>IN_0</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>8</ID>
<type>AM_REGISTER16</type>
<position>-6,-70.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>116 </input>
<input>
<ID>IN_10</ID>115 </input>
<input>
<ID>IN_11</ID>120 </input>
<input>
<ID>IN_12</ID>122 </input>
<input>
<ID>IN_13</ID>117 </input>
<input>
<ID>IN_14</ID>118 </input>
<input>
<ID>IN_15</ID>121 </input>
<input>
<ID>IN_2</ID>123 </input>
<input>
<ID>IN_3</ID>112 </input>
<input>
<ID>IN_4</ID>126 </input>
<input>
<ID>IN_5</ID>119 </input>
<input>
<ID>IN_6</ID>114 </input>
<input>
<ID>IN_7</ID>113 </input>
<input>
<ID>IN_8</ID>111 </input>
<input>
<ID>IN_9</ID>124 </input>
<output>
<ID>OUT_0</ID>369 </output>
<output>
<ID>OUT_1</ID>374 </output>
<output>
<ID>OUT_10</ID>377 </output>
<output>
<ID>OUT_11</ID>379 </output>
<output>
<ID>OUT_12</ID>380 </output>
<output>
<ID>OUT_13</ID>381 </output>
<output>
<ID>OUT_14</ID>371 </output>
<output>
<ID>OUT_15</ID>382 </output>
<output>
<ID>OUT_2</ID>375 </output>
<output>
<ID>OUT_3</ID>367 </output>
<output>
<ID>OUT_4</ID>373 </output>
<output>
<ID>OUT_5</ID>372 </output>
<output>
<ID>OUT_6</ID>368 </output>
<output>
<ID>OUT_7</ID>378 </output>
<output>
<ID>OUT_8</ID>370 </output>
<output>
<ID>OUT_9</ID>376 </output>
<input>
<ID>clear</ID>573 </input>
<input>
<ID>clock</ID>497 </input>
<input>
<ID>count_enable</ID>575 </input>
<input>
<ID>count_up</ID>574 </input>
<input>
<ID>load</ID>576 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>32.5,-39.5</position>
<gparam>LABEL_TEXT Program Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>-5.5,-54</position>
<gparam>LABEL_TEXT Data Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>31.5,-144.5</position>
<input>
<ID>IN_0</ID>494 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>36.5,-73.5</position>
<gparam>LABEL_TEXT Accumulator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>-10,-124.5</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>16</ID>
<type>AM_REGISTER16</type>
<position>-6.5,-111.5</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_10</ID>147 </input>
<input>
<ID>IN_11</ID>145 </input>
<input>
<ID>IN_12</ID>152 </input>
<input>
<ID>IN_13</ID>153 </input>
<input>
<ID>IN_14</ID>155 </input>
<input>
<ID>IN_15</ID>158 </input>
<input>
<ID>IN_2</ID>150 </input>
<input>
<ID>IN_3</ID>149 </input>
<input>
<ID>IN_4</ID>148 </input>
<input>
<ID>IN_5</ID>156 </input>
<input>
<ID>IN_6</ID>143 </input>
<input>
<ID>IN_7</ID>154 </input>
<input>
<ID>IN_8</ID>151 </input>
<input>
<ID>IN_9</ID>157 </input>
<output>
<ID>OUT_0</ID>431 </output>
<output>
<ID>OUT_1</ID>432 </output>
<output>
<ID>OUT_10</ID>439 </output>
<output>
<ID>OUT_11</ID>444 </output>
<output>
<ID>OUT_12</ID>443 </output>
<output>
<ID>OUT_13</ID>445 </output>
<output>
<ID>OUT_14</ID>442 </output>
<output>
<ID>OUT_15</ID>446 </output>
<output>
<ID>OUT_2</ID>433 </output>
<output>
<ID>OUT_3</ID>434 </output>
<output>
<ID>OUT_4</ID>435 </output>
<output>
<ID>OUT_5</ID>440 </output>
<output>
<ID>OUT_6</ID>441 </output>
<output>
<ID>OUT_7</ID>436 </output>
<output>
<ID>OUT_8</ID>437 </output>
<output>
<ID>OUT_9</ID>438 </output>
<input>
<ID>clock</ID>495 </input>
<input>
<ID>count_up</ID>579 </input>
<input>
<ID>load</ID>585 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>32,-102.5</position>
<input>
<ID>IN_0</ID>496 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>-6,-96.5</position>
<gparam>LABEL_TEXT Instruction Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>-10,-83</position>
<input>
<ID>IN_0</ID>497 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>18</ID>
<type>AM_REGISTER16</type>
<position>35.5,-131.5</position>
<input>
<ID>IN_0</ID>164 </input>
<input>
<ID>IN_1</ID>168 </input>
<input>
<ID>IN_10</ID>171 </input>
<input>
<ID>IN_11</ID>172 </input>
<input>
<ID>IN_12</ID>174 </input>
<input>
<ID>IN_13</ID>159 </input>
<input>
<ID>IN_14</ID>162 </input>
<input>
<ID>IN_15</ID>163 </input>
<input>
<ID>IN_2</ID>169 </input>
<input>
<ID>IN_3</ID>165 </input>
<input>
<ID>IN_4</ID>173 </input>
<input>
<ID>IN_5</ID>161 </input>
<input>
<ID>IN_6</ID>167 </input>
<input>
<ID>IN_7</ID>160 </input>
<input>
<ID>IN_8</ID>170 </input>
<input>
<ID>IN_9</ID>166 </input>
<output>
<ID>OUT_0</ID>465 </output>
<output>
<ID>OUT_1</ID>467 </output>
<output>
<ID>OUT_10</ID>469 </output>
<output>
<ID>OUT_11</ID>474 </output>
<output>
<ID>OUT_12</ID>478 </output>
<output>
<ID>OUT_13</ID>470 </output>
<output>
<ID>OUT_14</ID>472 </output>
<output>
<ID>OUT_15</ID>476 </output>
<output>
<ID>OUT_2</ID>463 </output>
<output>
<ID>OUT_3</ID>464 </output>
<output>
<ID>OUT_4</ID>466 </output>
<output>
<ID>OUT_5</ID>475 </output>
<output>
<ID>OUT_6</ID>477 </output>
<output>
<ID>OUT_7</ID>468 </output>
<output>
<ID>OUT_8</ID>471 </output>
<output>
<ID>OUT_9</ID>473 </output>
<input>
<ID>clear</ID>589 </input>
<input>
<ID>clock</ID>494 </input>
<input>
<ID>count_enable</ID>587 </input>
<input>
<ID>load</ID>588 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>36,-63</position>
<input>
<ID>IN_0</ID>498 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>36,-115</position>
<gparam>LABEL_TEXT Temporary Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>-5,-42</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>4,-136.5</position>
<gparam>LABEL_TEXT Output Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>BX_16X1_BUS_END</type>
<position>34.5,-29.5</position>
<input>
<ID>Bus_in_0</ID>294 </input>
<input>
<ID>IN_1</ID>293 </input>
<input>
<ID>IN_10</ID>282 </input>
<input>
<ID>IN_11</ID>281 </input>
<input>
<ID>IN_2</ID>292 </input>
<input>
<ID>IN_3</ID>291 </input>
<input>
<ID>IN_4</ID>290 </input>
<input>
<ID>IN_5</ID>289 </input>
<input>
<ID>IN_6</ID>288 </input>
<input>
<ID>IN_7</ID>287 </input>
<input>
<ID>IN_8</ID>279 </input>
<input>
<ID>IN_9</ID>280 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>25</ID>
<type>BX_16X1_BUS_END</type>
<position>23,-1</position>
<input>
<ID>Bus_in_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_10</ID>13 </input>
<input>
<ID>IN_11</ID>15 </input>
<input>
<ID>IN_12</ID>10 </input>
<input>
<ID>IN_13</ID>9 </input>
<input>
<ID>IN_14</ID>12 </input>
<input>
<ID>IN_15</ID>17 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>3 </input>
<input>
<ID>IN_4</ID>4 </input>
<input>
<ID>IN_5</ID>8 </input>
<input>
<ID>IN_6</ID>5 </input>
<input>
<ID>IN_7</ID>11 </input>
<input>
<ID>IN_8</ID>16 </input>
<input>
<ID>IN_9</ID>14 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>32</ID>
<type>BB_CLOCK</type>
<position>-19,4.5</position>
<output>
<ID>CLK</ID>492 </output>
<gparam>angle 0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>33</ID>
<type>BX_16X1_BUS_END</type>
<position>24.5,-51</position>
<input>
<ID>Bus_in_0</ID>108 </input>
<input>
<ID>IN_1</ID>107 </input>
<input>
<ID>IN_10</ID>106 </input>
<input>
<ID>IN_11</ID>101 </input>
<input>
<ID>IN_2</ID>109 </input>
<input>
<ID>IN_3</ID>110 </input>
<input>
<ID>IN_4</ID>99 </input>
<input>
<ID>IN_5</ID>104 </input>
<input>
<ID>IN_6</ID>105 </input>
<input>
<ID>IN_7</ID>100 </input>
<input>
<ID>IN_8</ID>103 </input>
<input>
<ID>IN_9</ID>102 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>34</ID>
<type>BX_16X1_BUS_END</type>
<position>-13.5,-70.5</position>
<input>
<ID>Bus_in_0</ID>125 </input>
<input>
<ID>IN_1</ID>116 </input>
<input>
<ID>IN_10</ID>115 </input>
<input>
<ID>IN_11</ID>120 </input>
<input>
<ID>IN_12</ID>122 </input>
<input>
<ID>IN_13</ID>117 </input>
<input>
<ID>IN_14</ID>118 </input>
<input>
<ID>IN_15</ID>121 </input>
<input>
<ID>IN_2</ID>123 </input>
<input>
<ID>IN_3</ID>112 </input>
<input>
<ID>IN_4</ID>126 </input>
<input>
<ID>IN_5</ID>119 </input>
<input>
<ID>IN_6</ID>114 </input>
<input>
<ID>IN_7</ID>113 </input>
<input>
<ID>IN_8</ID>111 </input>
<input>
<ID>IN_9</ID>124 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>99</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>48,-55</position>
<input>
<ID>ENABLE_0</ID>693 </input>
<input>
<ID>IN_0</ID>552 </input>
<input>
<ID>IN_1</ID>557 </input>
<input>
<ID>IN_2</ID>551 </input>
<input>
<ID>IN_3</ID>556 </input>
<input>
<ID>IN_4</ID>553 </input>
<input>
<ID>IN_5</ID>554 </input>
<input>
<ID>IN_6</ID>555 </input>
<input>
<ID>IN_7</ID>558 </input>
<output>
<ID>OUT_0</ID>661 </output>
<output>
<ID>OUT_1</ID>662 </output>
<output>
<ID>OUT_2</ID>663 </output>
<output>
<ID>OUT_3</ID>664 </output>
<output>
<ID>OUT_4</ID>665 </output>
<output>
<ID>OUT_5</ID>666 </output>
<output>
<ID>OUT_6</ID>667 </output>
<output>
<ID>OUT_7</ID>668 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>36</ID>
<type>BX_16X1_BUS_END</type>
<position>-14,-111.5</position>
<input>
<ID>Bus_in_0</ID>146 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_10</ID>147 </input>
<input>
<ID>IN_11</ID>145 </input>
<input>
<ID>IN_12</ID>152 </input>
<input>
<ID>IN_13</ID>153 </input>
<input>
<ID>IN_14</ID>155 </input>
<input>
<ID>IN_15</ID>158 </input>
<input>
<ID>IN_2</ID>150 </input>
<input>
<ID>IN_3</ID>149 </input>
<input>
<ID>IN_4</ID>148 </input>
<input>
<ID>IN_5</ID>156 </input>
<input>
<ID>IN_6</ID>143 </input>
<input>
<ID>IN_7</ID>154 </input>
<input>
<ID>IN_8</ID>151 </input>
<input>
<ID>IN_9</ID>157 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>100</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>52.5,-49</position>
<input>
<ID>ENABLE_0</ID>693 </input>
<input>
<ID>IN_0</ID>559 </input>
<input>
<ID>IN_1</ID>560 </input>
<input>
<ID>IN_2</ID>561 </input>
<input>
<ID>IN_3</ID>562 </input>
<output>
<ID>OUT_0</ID>657 </output>
<output>
<ID>OUT_1</ID>658 </output>
<output>
<ID>OUT_2</ID>660 </output>
<output>
<ID>OUT_3</ID>659 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>37</ID>
<type>BX_16X1_BUS_END</type>
<position>28,-131.5</position>
<input>
<ID>Bus_in_0</ID>164 </input>
<input>
<ID>IN_1</ID>168 </input>
<input>
<ID>IN_10</ID>171 </input>
<input>
<ID>IN_11</ID>172 </input>
<input>
<ID>IN_12</ID>174 </input>
<input>
<ID>IN_13</ID>159 </input>
<input>
<ID>IN_14</ID>162 </input>
<input>
<ID>IN_15</ID>163 </input>
<input>
<ID>IN_2</ID>169 </input>
<input>
<ID>IN_3</ID>165 </input>
<input>
<ID>IN_4</ID>173 </input>
<input>
<ID>IN_5</ID>161 </input>
<input>
<ID>IN_6</ID>167 </input>
<input>
<ID>IN_7</ID>160 </input>
<input>
<ID>IN_8</ID>170 </input>
<input>
<ID>IN_9</ID>166 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>117</ID>
<type>DA_FROM</type>
<position>-3,-57.5</position>
<input>
<ID>IN_0</ID>575 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID inc_dr</lparam></gate>
<gate>
<ID>53</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>1.5,-70.5</position>
<input>
<ID>ENABLE_0</ID>694 </input>
<input>
<ID>IN_0</ID>369 </input>
<input>
<ID>IN_1</ID>374 </input>
<input>
<ID>IN_10</ID>377 </input>
<input>
<ID>IN_11</ID>379 </input>
<input>
<ID>IN_12</ID>380 </input>
<input>
<ID>IN_13</ID>381 </input>
<input>
<ID>IN_14</ID>371 </input>
<input>
<ID>IN_15</ID>382 </input>
<input>
<ID>IN_2</ID>375 </input>
<input>
<ID>IN_3</ID>367 </input>
<input>
<ID>IN_4</ID>373 </input>
<input>
<ID>IN_5</ID>372 </input>
<input>
<ID>IN_6</ID>368 </input>
<input>
<ID>IN_7</ID>378 </input>
<input>
<ID>IN_8</ID>370 </input>
<input>
<ID>IN_9</ID>376 </input>
<output>
<ID>OUT_0</ID>365 </output>
<output>
<ID>OUT_1</ID>366 </output>
<output>
<ID>OUT_10</ID>352 </output>
<output>
<ID>OUT_11</ID>357 </output>
<output>
<ID>OUT_12</ID>351 </output>
<output>
<ID>OUT_13</ID>358 </output>
<output>
<ID>OUT_14</ID>356 </output>
<output>
<ID>OUT_15</ID>359 </output>
<output>
<ID>OUT_2</ID>362 </output>
<output>
<ID>OUT_3</ID>363 </output>
<output>
<ID>OUT_4</ID>360 </output>
<output>
<ID>OUT_5</ID>361 </output>
<output>
<ID>OUT_6</ID>364 </output>
<output>
<ID>OUT_7</ID>353 </output>
<output>
<ID>OUT_8</ID>354 </output>
<output>
<ID>OUT_9</ID>355 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>118</ID>
<type>EE_VDD</type>
<position>-5,-59.5</position>
<output>
<ID>OUT_0</ID>574 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>54</ID>
<type>BX_16X1_BUS_END</type>
<position>6,-70.5</position>
<input>
<ID>Bus_in_0</ID>365 </input>
<input>
<ID>IN_1</ID>366 </input>
<input>
<ID>IN_10</ID>352 </input>
<input>
<ID>IN_11</ID>357 </input>
<input>
<ID>IN_12</ID>351 </input>
<input>
<ID>IN_13</ID>358 </input>
<input>
<ID>IN_14</ID>356 </input>
<input>
<ID>IN_15</ID>359 </input>
<input>
<ID>IN_2</ID>362 </input>
<input>
<ID>IN_3</ID>363 </input>
<input>
<ID>IN_4</ID>360 </input>
<input>
<ID>IN_5</ID>361 </input>
<input>
<ID>IN_6</ID>364 </input>
<input>
<ID>IN_7</ID>353 </input>
<input>
<ID>IN_8</ID>354 </input>
<input>
<ID>IN_9</ID>355 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>119</ID>
<type>DA_FROM</type>
<position>-10.5,-59.5</position>
<input>
<ID>IN_0</ID>576 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_dr</lparam></gate>
<gate>
<ID>55</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>43.5,-90</position>
<input>
<ID>ENABLE_0</ID>695 </input>
<input>
<ID>IN_0</ID>414 </input>
<input>
<ID>IN_1</ID>399 </input>
<input>
<ID>IN_10</ID>405 </input>
<input>
<ID>IN_11</ID>403 </input>
<input>
<ID>IN_12</ID>404 </input>
<input>
<ID>IN_13</ID>406 </input>
<input>
<ID>IN_14</ID>407 </input>
<input>
<ID>IN_15</ID>409 </input>
<input>
<ID>IN_2</ID>410 </input>
<input>
<ID>IN_3</ID>400 </input>
<input>
<ID>IN_4</ID>401 </input>
<input>
<ID>IN_5</ID>408 </input>
<input>
<ID>IN_6</ID>411 </input>
<input>
<ID>IN_7</ID>412 </input>
<input>
<ID>IN_8</ID>402 </input>
<input>
<ID>IN_9</ID>413 </input>
<output>
<ID>OUT_0</ID>397 </output>
<output>
<ID>OUT_1</ID>398 </output>
<output>
<ID>OUT_10</ID>384 </output>
<output>
<ID>OUT_11</ID>389 </output>
<output>
<ID>OUT_12</ID>383 </output>
<output>
<ID>OUT_13</ID>390 </output>
<output>
<ID>OUT_14</ID>388 </output>
<output>
<ID>OUT_15</ID>391 </output>
<output>
<ID>OUT_2</ID>394 </output>
<output>
<ID>OUT_3</ID>395 </output>
<output>
<ID>OUT_4</ID>392 </output>
<output>
<ID>OUT_5</ID>393 </output>
<output>
<ID>OUT_6</ID>396 </output>
<output>
<ID>OUT_7</ID>385 </output>
<output>
<ID>OUT_8</ID>386 </output>
<output>
<ID>OUT_9</ID>387 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>120</ID>
<type>DA_FROM</type>
<position>38.5,-77</position>
<input>
<ID>IN_0</ID>577 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID inc_ac</lparam></gate>
<gate>
<ID>56</ID>
<type>BX_16X1_BUS_END</type>
<position>48,-90</position>
<input>
<ID>Bus_in_0</ID>397 </input>
<input>
<ID>IN_1</ID>398 </input>
<input>
<ID>IN_10</ID>384 </input>
<input>
<ID>IN_11</ID>389 </input>
<input>
<ID>IN_12</ID>383 </input>
<input>
<ID>IN_13</ID>390 </input>
<input>
<ID>IN_14</ID>388 </input>
<input>
<ID>IN_15</ID>391 </input>
<input>
<ID>IN_2</ID>394 </input>
<input>
<ID>IN_3</ID>395 </input>
<input>
<ID>IN_4</ID>392 </input>
<input>
<ID>IN_5</ID>393 </input>
<input>
<ID>IN_6</ID>396 </input>
<input>
<ID>IN_7</ID>385 </input>
<input>
<ID>IN_8</ID>386 </input>
<input>
<ID>IN_9</ID>387 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>121</ID>
<type>EE_VDD</type>
<position>37,-79</position>
<output>
<ID>OUT_0</ID>578 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>57</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>1,-111.5</position>
<input>
<ID>ENABLE_0</ID>696 </input>
<input>
<ID>IN_0</ID>431 </input>
<input>
<ID>IN_1</ID>432 </input>
<input>
<ID>IN_10</ID>439 </input>
<input>
<ID>IN_11</ID>444 </input>
<input>
<ID>IN_12</ID>443 </input>
<input>
<ID>IN_13</ID>445 </input>
<input>
<ID>IN_14</ID>442 </input>
<input>
<ID>IN_15</ID>446 </input>
<input>
<ID>IN_2</ID>433 </input>
<input>
<ID>IN_3</ID>434 </input>
<input>
<ID>IN_4</ID>435 </input>
<input>
<ID>IN_5</ID>440 </input>
<input>
<ID>IN_6</ID>441 </input>
<input>
<ID>IN_7</ID>436 </input>
<input>
<ID>IN_8</ID>437 </input>
<input>
<ID>IN_9</ID>438 </input>
<output>
<ID>OUT_0</ID>429 </output>
<output>
<ID>OUT_1</ID>430 </output>
<output>
<ID>OUT_10</ID>416 </output>
<output>
<ID>OUT_11</ID>421 </output>
<output>
<ID>OUT_12</ID>415 </output>
<output>
<ID>OUT_13</ID>422 </output>
<output>
<ID>OUT_14</ID>420 </output>
<output>
<ID>OUT_15</ID>423 </output>
<output>
<ID>OUT_2</ID>426 </output>
<output>
<ID>OUT_3</ID>427 </output>
<output>
<ID>OUT_4</ID>424 </output>
<output>
<ID>OUT_5</ID>425 </output>
<output>
<ID>OUT_6</ID>428 </output>
<output>
<ID>OUT_8</ID>418 </output>
<output>
<ID>OUT_9</ID>419 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>122</ID>
<type>EE_VDD</type>
<position>-5.5,-100.5</position>
<output>
<ID>OUT_0</ID>579 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>58</ID>
<type>BX_16X1_BUS_END</type>
<position>5.5,-111.5</position>
<input>
<ID>Bus_in_0</ID>429 </input>
<input>
<ID>IN_1</ID>430 </input>
<input>
<ID>IN_10</ID>416 </input>
<input>
<ID>IN_11</ID>421 </input>
<input>
<ID>IN_12</ID>415 </input>
<input>
<ID>IN_13</ID>422 </input>
<input>
<ID>IN_14</ID>420 </input>
<input>
<ID>IN_15</ID>423 </input>
<input>
<ID>IN_2</ID>426 </input>
<input>
<ID>IN_3</ID>427 </input>
<input>
<ID>IN_4</ID>424 </input>
<input>
<ID>IN_5</ID>425 </input>
<input>
<ID>IN_6</ID>428 </input>
<input>
<ID>IN_7</ID>417 </input>
<input>
<ID>IN_8</ID>418 </input>
<input>
<ID>IN_9</ID>419 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>59</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>43,-131.5</position>
<input>
<ID>ENABLE_0</ID>697 </input>
<input>
<ID>IN_0</ID>465 </input>
<input>
<ID>IN_1</ID>467 </input>
<input>
<ID>IN_10</ID>469 </input>
<input>
<ID>IN_11</ID>474 </input>
<input>
<ID>IN_12</ID>478 </input>
<input>
<ID>IN_13</ID>470 </input>
<input>
<ID>IN_14</ID>472 </input>
<input>
<ID>IN_15</ID>476 </input>
<input>
<ID>IN_2</ID>463 </input>
<input>
<ID>IN_3</ID>464 </input>
<input>
<ID>IN_4</ID>466 </input>
<input>
<ID>IN_5</ID>475 </input>
<input>
<ID>IN_6</ID>477 </input>
<input>
<ID>IN_7</ID>468 </input>
<input>
<ID>IN_8</ID>471 </input>
<input>
<ID>IN_9</ID>473 </input>
<output>
<ID>OUT_0</ID>461 </output>
<output>
<ID>OUT_1</ID>462 </output>
<output>
<ID>OUT_10</ID>448 </output>
<output>
<ID>OUT_11</ID>453 </output>
<output>
<ID>OUT_12</ID>447 </output>
<output>
<ID>OUT_13</ID>454 </output>
<output>
<ID>OUT_14</ID>452 </output>
<output>
<ID>OUT_15</ID>455 </output>
<output>
<ID>OUT_2</ID>458 </output>
<output>
<ID>OUT_3</ID>459 </output>
<output>
<ID>OUT_4</ID>456 </output>
<output>
<ID>OUT_5</ID>457 </output>
<output>
<ID>OUT_6</ID>460 </output>
<output>
<ID>OUT_7</ID>449 </output>
<output>
<ID>OUT_8</ID>450 </output>
<output>
<ID>OUT_9</ID>451 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>124</ID>
<type>EE_VDD</type>
<position>4.5,-141</position>
<output>
<ID>OUT_0</ID>581 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>60</ID>
<type>BX_16X1_BUS_END</type>
<position>47.5,-131.5</position>
<input>
<ID>Bus_in_0</ID>461 </input>
<input>
<ID>IN_1</ID>462 </input>
<input>
<ID>IN_10</ID>448 </input>
<input>
<ID>IN_11</ID>453 </input>
<input>
<ID>IN_12</ID>447 </input>
<input>
<ID>IN_13</ID>454 </input>
<input>
<ID>IN_14</ID>452 </input>
<input>
<ID>IN_15</ID>455 </input>
<input>
<ID>IN_2</ID>458 </input>
<input>
<ID>IN_3</ID>459 </input>
<input>
<ID>IN_4</ID>456 </input>
<input>
<ID>IN_5</ID>457 </input>
<input>
<ID>IN_6</ID>460 </input>
<input>
<ID>IN_7</ID>449 </input>
<input>
<ID>IN_8</ID>450 </input>
<input>
<ID>IN_9</ID>451 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>105</ID>
<type>DA_FROM</type>
<position>44.5,13</position>
<input>
<ID>IN_0</ID>563 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID mem_w</lparam></gate>
<gate>
<ID>106</ID>
<type>DA_FROM</type>
<position>34.5,12</position>
<input>
<ID>IN_0</ID>564 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID mem_r</lparam></gate>
<gate>
<ID>107</ID>
<type>DA_FROM</type>
<position>3,-42</position>
<input>
<ID>IN_0</ID>565 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clr_addr</lparam></gate>
<gate>
<ID>108</ID>
<type>DA_FROM</type>
<position>-4.5,-22.5</position>
<input>
<ID>IN_0</ID>566 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_addr</lparam></gate>
<gate>
<ID>111</ID>
<type>DA_FROM</type>
<position>2,-20.5</position>
<input>
<ID>IN_0</ID>568 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID inc_addr</lparam></gate>
<gate>
<ID>112</ID>
<type>DA_FROM</type>
<position>44,-63</position>
<input>
<ID>IN_0</ID>569 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clr_pc</lparam></gate>
<gate>
<ID>113</ID>
<type>DA_FROM</type>
<position>35,-44</position>
<input>
<ID>IN_0</ID>570 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_pc</lparam></gate>
<gate>
<ID>114</ID>
<type>DA_FROM</type>
<position>44,-43</position>
<input>
<ID>IN_0</ID>572 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID inc_pc</lparam></gate>
<gate>
<ID>115</ID>
<type>EE_VDD</type>
<position>41,-44</position>
<output>
<ID>OUT_0</ID>571 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>116</ID>
<type>DA_FROM</type>
<position>-2,-83</position>
<input>
<ID>IN_0</ID>573 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clr_data</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>31,-79</position>
<input>
<ID>IN_0</ID>582 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_ac</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>40,-102.5</position>
<input>
<ID>IN_0</ID>583 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clr_ac</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>-10.5,-101</position>
<input>
<ID>IN_0</ID>585 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_ir</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>31,-120.5</position>
<input>
<ID>IN_0</ID>588 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_tr</lparam></gate>
<gate>
<ID>136</ID>
<type>BX_16X1_BUS_END</type>
<position>-11.5,-144</position>
<input>
<ID>Bus_in_0</ID>609 </input>
<input>
<ID>IN_1</ID>610 </input>
<input>
<ID>IN_2</ID>611 </input>
<input>
<ID>IN_3</ID>614 </input>
<input>
<ID>IN_4</ID>615 </input>
<input>
<ID>IN_5</ID>616 </input>
<input>
<ID>IN_6</ID>612 </input>
<input>
<ID>IN_7</ID>613 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>137</ID>
<type>BX_16X1_BUS_END</type>
<position>61.5,-51</position>
<input>
<ID>Bus_in_0</ID>661 </input>
<input>
<ID>IN_1</ID>662 </input>
<input>
<ID>IN_10</ID>660 </input>
<input>
<ID>IN_11</ID>659 </input>
<input>
<ID>IN_2</ID>663 </input>
<input>
<ID>IN_3</ID>664 </input>
<input>
<ID>IN_4</ID>665 </input>
<input>
<ID>IN_5</ID>666 </input>
<input>
<ID>IN_6</ID>667 </input>
<input>
<ID>IN_7</ID>668 </input>
<input>
<ID>IN_8</ID>657 </input>
<input>
<ID>IN_9</ID>658 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>164</ID>
<type>DA_FROM</type>
<position>55.5,-40</position>
<input>
<ID>IN_0</ID>693 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_pc</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>8,-59.5</position>
<input>
<ID>IN_0</ID>694 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_dr</lparam></gate>
<gate>
<ID>166</ID>
<type>DA_FROM</type>
<position>51.5,-79</position>
<input>
<ID>IN_0</ID>695 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_ac</lparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>7,-100.5</position>
<input>
<ID>IN_0</ID>696 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_ir</lparam></gate>
<gate>
<ID>168</ID>
<type>DA_FROM</type>
<position>48,-119.5</position>
<input>
<ID>IN_0</ID>697 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_tr</lparam></gate>
<gate>
<ID>27</ID>
<type>BX_16X1_BUS_END</type>
<position>-15.5,-29.5</position>
<input>
<ID>Bus_in_0</ID>95 </input>
<input>
<ID>IN_1</ID>179 </input>
<input>
<ID>IN_10</ID>177 </input>
<input>
<ID>IN_11</ID>178 </input>
<input>
<ID>IN_2</ID>93 </input>
<input>
<ID>IN_3</ID>96 </input>
<input>
<ID>IN_4</ID>97 </input>
<input>
<ID>IN_5</ID>98 </input>
<input>
<ID>IN_6</ID>176 </input>
<input>
<ID>IN_7</ID>94 </input>
<input>
<ID>IN_8</ID>180 </input>
<input>
<ID>IN_9</ID>175 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>66</ID>
<type>BX_16X1_BUS_END</type>
<position>9,-29.5</position>
<input>
<ID>Bus_in_0</ID>188 </input>
<input>
<ID>IN_1</ID>182 </input>
<input>
<ID>IN_10</ID>191 </input>
<input>
<ID>IN_11</ID>192 </input>
<input>
<ID>IN_2</ID>190 </input>
<input>
<ID>IN_3</ID>189 </input>
<input>
<ID>IN_4</ID>181 </input>
<input>
<ID>IN_5</ID>183 </input>
<input>
<ID>IN_6</ID>184 </input>
<input>
<ID>IN_7</ID>185 </input>
<input>
<ID>IN_8</ID>187 </input>
<input>
<ID>IN_9</ID>186 </input>
<input>
<ID>OUT</ID>205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>67</ID>
<type>BX_16X1_BUS_END</type>
<position>10.5,14.5</position>
<input>
<ID>Bus_in_0</ID>197 </input>
<input>
<ID>IN_1</ID>198 </input>
<input>
<ID>IN_10</ID>203 </input>
<input>
<ID>IN_11</ID>204 </input>
<input>
<ID>IN_2</ID>195 </input>
<input>
<ID>IN_3</ID>201 </input>
<input>
<ID>IN_4</ID>199 </input>
<input>
<ID>IN_5</ID>202 </input>
<input>
<ID>IN_6</ID>200 </input>
<input>
<ID>IN_7</ID>193 </input>
<input>
<ID>IN_8</ID>194 </input>
<input>
<ID>IN_9</ID>196 </input>
<input>
<ID>OUT</ID>205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>68</ID>
<type>BX_16X1_BUS_END</type>
<position>20.5,-29.5</position>
<input>
<ID>Bus_in_0</ID>272 </input>
<input>
<ID>IN_1</ID>276 </input>
<input>
<ID>IN_10</ID>285 </input>
<input>
<ID>IN_11</ID>286 </input>
<input>
<ID>IN_2</ID>273 </input>
<input>
<ID>IN_3</ID>275 </input>
<input>
<ID>IN_4</ID>277 </input>
<input>
<ID>IN_5</ID>271 </input>
<input>
<ID>IN_6</ID>274 </input>
<input>
<ID>IN_7</ID>278 </input>
<input>
<ID>IN_8</ID>283 </input>
<input>
<ID>IN_9</ID>284 </input>
<input>
<ID>OUT</ID>205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>33,-18</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_ar</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>28.5,-97.5</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc0</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>19.5,-96.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc1</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>28.5,-95.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc2</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>19.5,-94.5</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc3</lparam></gate>
<gate>
<ID>85</ID>
<type>DA_FROM</type>
<position>28.5,-93.5</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc4</lparam></gate>
<gate>
<ID>86</ID>
<type>DA_FROM</type>
<position>19.5,-92.5</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc5</lparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>28.5,-91.5</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc6</lparam></gate>
<gate>
<ID>88</ID>
<type>DA_FROM</type>
<position>19.5,-90.5</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc7</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>28.5,-89.5</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc8</lparam></gate>
<gate>
<ID>90</ID>
<type>DA_FROM</type>
<position>19.5,-88.5</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc9</lparam></gate>
<gate>
<ID>91</ID>
<type>DA_FROM</type>
<position>28.5,-87.5</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc10</lparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>19.5,-86.5</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc11</lparam></gate>
<gate>
<ID>93</ID>
<type>DA_FROM</type>
<position>28.5,-85.5</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc12</lparam></gate>
<gate>
<ID>94</ID>
<type>DA_FROM</type>
<position>19.5,-84.5</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc13</lparam></gate>
<gate>
<ID>95</ID>
<type>DA_FROM</type>
<position>28.5,-83.5</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc14</lparam></gate>
<gate>
<ID>96</ID>
<type>DA_FROM</type>
<position>19.5,-82.5</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc15</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>-60.5,20.5</position>
<gparam>LABEL_TEXT Mano Machine</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>-52,14</position>
<gparam>LABEL_TEXT Checkpoint 1 - Brandon Aikman</gparam>
<gparam>TEXT_HEIGHT 2.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>25.5,-33.5</position>
<input>
<ID>ENABLE_0</ID>295 </input>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>276 </input>
<input>
<ID>IN_2</ID>273 </input>
<input>
<ID>IN_3</ID>275 </input>
<input>
<ID>IN_4</ID>277 </input>
<input>
<ID>IN_5</ID>271 </input>
<input>
<ID>IN_6</ID>274 </input>
<input>
<ID>IN_7</ID>278 </input>
<output>
<ID>OUT_0</ID>294 </output>
<output>
<ID>OUT_1</ID>293 </output>
<output>
<ID>OUT_2</ID>292 </output>
<output>
<ID>OUT_3</ID>291 </output>
<output>
<ID>OUT_4</ID>290 </output>
<output>
<ID>OUT_5</ID>289 </output>
<output>
<ID>OUT_6</ID>288 </output>
<output>
<ID>OUT_7</ID>287 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>102</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>30,-27.5</position>
<input>
<ID>ENABLE_0</ID>295 </input>
<input>
<ID>IN_0</ID>283 </input>
<input>
<ID>IN_1</ID>284 </input>
<input>
<ID>IN_2</ID>285 </input>
<input>
<ID>IN_3</ID>286 </input>
<output>
<ID>OUT_0</ID>279 </output>
<output>
<ID>OUT_1</ID>280 </output>
<output>
<ID>OUT_2</ID>282 </output>
<output>
<ID>OUT_3</ID>281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>414 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-97.5,41.5,-97.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>563 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,13,42.5,13</points>
<connection>
<GID>2</GID>
<name>write_enable</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,1,24.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_6</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>25</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>197 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,7,14,7</points>
<connection>
<GID>2</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>67</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>572 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-45.5,40,-43</points>
<connection>
<GID>12</GID>
<name>count_enable</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-43,42,-43</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>6 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,1,30.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_0</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>Bus_in_0</name></connection></vsegment></shape></wire>
<wire>
<ID>493 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-158,2.5,-153.5</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<intersection>-158 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-158,2.5,-158</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>198 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,8,14,8</points>
<connection>
<GID>2</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>67</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>3 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,1,27.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_3</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>25</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>356 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-64,4,-64</points>
<connection>
<GID>53</GID>
<name>OUT_14</name></connection>
<connection>
<GID>54</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>195 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,9,14,9</points>
<connection>
<GID>2</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>67</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>492 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-15,4.5,-9,4.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>11 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,1,23.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_7</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>25</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>364 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-72,4,-72</points>
<connection>
<GID>53</GID>
<name>OUT_6</name></connection>
<connection>
<GID>54</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>203 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,17,14,17</points>
<connection>
<GID>2</GID>
<name>ADDRESS_10</name></connection>
<connection>
<GID>67</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>12 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,1,16.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_14</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_14</name></connection>
<connection>
<GID>25</GID>
<name>IN_14</name></connection></vsegment></shape></wire>
<wire>
<ID>491 </ID>
<shape>
<hsegment>
<ID>8</ID>
<points>32,14,32.5,14</points>
<connection>
<GID>2</GID>
<name>write_clock</name></connection>
<connection>
<GID>74</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>204 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,18,14,18</points>
<connection>
<GID>2</GID>
<name>ADDRESS_11</name></connection>
<connection>
<GID>67</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>9 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,1,17.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_13</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_13</name></connection>
<connection>
<GID>25</GID>
<name>IN_13</name></connection></vsegment></shape></wire>
<wire>
<ID>354 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-70,4,-70</points>
<connection>
<GID>53</GID>
<name>OUT_8</name></connection>
<connection>
<GID>54</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>201 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,10,14,10</points>
<connection>
<GID>2</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>67</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>7 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,1,29.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_1</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>25</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>199 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,11,14,11</points>
<connection>
<GID>2</GID>
<name>ADDRESS_4</name></connection>
<connection>
<GID>67</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>497 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-83,-7,-80</points>
<connection>
<GID>8</GID>
<name>clock</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,-83,-7,-83</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>10 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,1,18.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_12</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_12</name></connection>
<connection>
<GID>25</GID>
<name>IN_12</name></connection></vsegment></shape></wire>
<wire>
<ID>202 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,12,14,12</points>
<connection>
<GID>2</GID>
<name>ADDRESS_5</name></connection>
<connection>
<GID>67</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>8 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,1,25.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_5</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>25</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>200 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,13,14,13</points>
<connection>
<GID>2</GID>
<name>ADDRESS_6</name></connection>
<connection>
<GID>67</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>193 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,14,14,14</points>
<connection>
<GID>2</GID>
<name>ADDRESS_7</name></connection>
<connection>
<GID>67</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>2 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,1,28.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_2</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>25</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>194 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,15,14,15</points>
<connection>
<GID>2</GID>
<name>ADDRESS_8</name></connection>
<connection>
<GID>67</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>4 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,1,26.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_4</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>25</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>196 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,16,14,16</points>
<connection>
<GID>2</GID>
<name>ADDRESS_9</name></connection>
<connection>
<GID>67</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>422 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-106,3.5,-106</points>
<connection>
<GID>57</GID>
<name>OUT_13</name></connection>
<connection>
<GID>58</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>571 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-45.5,41,-45</points>
<connection>
<GID>12</GID>
<name>count_up</name></connection>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,1,20.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_10</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_10</name></connection>
<connection>
<GID>25</GID>
<name>IN_10</name></connection></vsegment></shape></wire>
<wire>
<ID>15 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,1,19.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_11</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_11</name></connection>
<connection>
<GID>25</GID>
<name>IN_11</name></connection></vsegment></shape></wire>
<wire>
<ID>591 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-142.5,2.5,-141</points>
<connection>
<GID>4</GID>
<name>load</name></connection>
<intersection>-141 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-141,2.5,-141</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,1,15.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_15</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_15</name></connection>
<connection>
<GID>25</GID>
<name>IN_15</name></connection></vsegment></shape></wire>
<wire>
<ID>16 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,1,22.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_8</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_8</name></connection>
<connection>
<GID>25</GID>
<name>IN_8</name></connection></vsegment></shape></wire>
<wire>
<ID>14 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,1,21.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_9</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_9</name></connection>
<connection>
<GID>25</GID>
<name>IN_9</name></connection></vsegment></shape></wire>
<wire>
<ID>564 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,12,32.5,12</points>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>432 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-118,-1,-118</points>
<connection>
<GID>16</GID>
<name>OUT_1</name></connection>
<connection>
<GID>57</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>609 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-151.5,-0.5,-151.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>136</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>610 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-150.5,-0.5,-150.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>136</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>462 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-138,45.5,-138</points>
<connection>
<GID>59</GID>
<name>OUT_1</name></connection>
<connection>
<GID>60</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>611 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-149.5,-0.5,-149.5</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<connection>
<GID>136</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>614 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-148.5,-0.5,-148.5</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<connection>
<GID>136</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>386 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-89.5,46,-89.5</points>
<connection>
<GID>55</GID>
<name>OUT_8</name></connection>
<connection>
<GID>56</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>551 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-56.5,46,-56.5</points>
<connection>
<GID>12</GID>
<name>OUT_2</name></connection>
<connection>
<GID>99</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>105 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-52.5,35,-52.5</points>
<connection>
<GID>12</GID>
<name>IN_6</name></connection>
<connection>
<GID>33</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>450 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-131,45.5,-131</points>
<connection>
<GID>59</GID>
<name>OUT_8</name></connection>
<connection>
<GID>60</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>615 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-147.5,-0.5,-147.5</points>
<connection>
<GID>4</GID>
<name>IN_4</name></connection>
<connection>
<GID>136</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>552 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-58.5,46,-58.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>281 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32,-26,32.5,-26</points>
<connection>
<GID>102</GID>
<name>OUT_3</name></connection>
<connection>
<GID>24</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>616 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-146.5,-0.5,-146.5</points>
<connection>
<GID>4</GID>
<name>IN_5</name></connection>
<connection>
<GID>136</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>469 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-129,41,-129</points>
<connection>
<GID>18</GID>
<name>OUT_10</name></connection>
<connection>
<GID>59</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>110 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-55.5,35,-55.5</points>
<connection>
<GID>12</GID>
<name>IN_3</name></connection>
<connection>
<GID>33</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>277 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-33,23.5,-33</points>
<connection>
<GID>68</GID>
<name>IN_4</name></connection>
<connection>
<GID>101</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>612 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-145.5,-0.5,-145.5</points>
<connection>
<GID>4</GID>
<name>IN_6</name></connection>
<connection>
<GID>136</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>436 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-112,-1,-112</points>
<connection>
<GID>16</GID>
<name>OUT_7</name></connection>
<connection>
<GID>57</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>613 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-144.5,-0.5,-144.5</points>
<connection>
<GID>4</GID>
<name>IN_7</name></connection>
<connection>
<GID>136</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>404 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-85.5,41.5,-85.5</points>
<connection>
<GID>14</GID>
<name>OUT_12</name></connection>
<connection>
<GID>55</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>581 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-142.5,4.5,-142</points>
<connection>
<GID>4</GID>
<name>count_up</name></connection>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>459 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-136,45.5,-136</points>
<connection>
<GID>59</GID>
<name>OUT_3</name></connection>
<connection>
<GID>60</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>108 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-58.5,35,-58.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>33</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>107 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-57.5,35,-57.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<connection>
<GID>33</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>465 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-139,41,-139</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>106 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-48.5,35,-48.5</points>
<connection>
<GID>12</GID>
<name>IN_10</name></connection>
<connection>
<GID>33</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>101 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-47.5,35,-47.5</points>
<connection>
<GID>12</GID>
<name>IN_11</name></connection>
<connection>
<GID>33</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>109 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-56.5,35,-56.5</points>
<connection>
<GID>12</GID>
<name>IN_2</name></connection>
<connection>
<GID>33</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>99 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-54.5,35,-54.5</points>
<connection>
<GID>12</GID>
<name>IN_4</name></connection>
<connection>
<GID>33</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>562 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-47.5,50.5,-47.5</points>
<connection>
<GID>12</GID>
<name>OUT_11</name></connection>
<connection>
<GID>100</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>471 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-131,41,-131</points>
<connection>
<GID>18</GID>
<name>OUT_8</name></connection>
<connection>
<GID>59</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>104 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-53.5,35,-53.5</points>
<connection>
<GID>12</GID>
<name>IN_5</name></connection>
<connection>
<GID>33</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>451 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-130,45.5,-130</points>
<connection>
<GID>59</GID>
<name>OUT_9</name></connection>
<connection>
<GID>60</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>100 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-51.5,35,-51.5</points>
<connection>
<GID>12</GID>
<name>IN_7</name></connection>
<connection>
<GID>33</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>103 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-50.5,35,-50.5</points>
<connection>
<GID>12</GID>
<name>IN_8</name></connection>
<connection>
<GID>33</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>461 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-139,45.5,-139</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<connection>
<GID>60</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>102 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-49.5,35,-49.5</points>
<connection>
<GID>12</GID>
<name>IN_9</name></connection>
<connection>
<GID>33</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>264 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-82.5,31,-82.5</points>
<connection>
<GID>14</GID>
<name>IN_15</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>569 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-63,41,-60.5</points>
<connection>
<GID>12</GID>
<name>clear</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-63,42,-63</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>498 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-63,39,-60.5</points>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-63,39,-63</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>570 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-45.5,39,-44</points>
<connection>
<GID>12</GID>
<name>load</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-44,39,-44</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>380 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-66,-0.5,-66</points>
<connection>
<GID>8</GID>
<name>OUT_12</name></connection>
<connection>
<GID>53</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>557 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-57.5,46,-57.5</points>
<connection>
<GID>12</GID>
<name>OUT_1</name></connection>
<connection>
<GID>99</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>256 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-95.5,31,-95.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<connection>
<GID>75</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>561 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-48.5,50.5,-48.5</points>
<connection>
<GID>12</GID>
<name>OUT_10</name></connection>
<connection>
<GID>100</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>556 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-55.5,46,-55.5</points>
<connection>
<GID>12</GID>
<name>OUT_3</name></connection>
<connection>
<GID>99</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>376 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-69,-0.5,-69</points>
<connection>
<GID>8</GID>
<name>OUT_9</name></connection>
<connection>
<GID>53</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>553 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-54.5,46,-54.5</points>
<connection>
<GID>12</GID>
<name>OUT_4</name></connection>
<connection>
<GID>99</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>554 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-53.5,46,-53.5</points>
<connection>
<GID>12</GID>
<name>OUT_5</name></connection>
<connection>
<GID>99</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>406 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-84.5,41.5,-84.5</points>
<connection>
<GID>14</GID>
<name>OUT_13</name></connection>
<connection>
<GID>55</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>555 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-52.5,46,-52.5</points>
<connection>
<GID>12</GID>
<name>OUT_6</name></connection>
<connection>
<GID>99</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>558 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-51.5,46,-51.5</points>
<connection>
<GID>12</GID>
<name>OUT_7</name></connection>
<connection>
<GID>99</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>394 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-95.5,46,-95.5</points>
<connection>
<GID>55</GID>
<name>OUT_2</name></connection>
<connection>
<GID>56</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>559 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-50.5,50.5,-50.5</points>
<connection>
<GID>12</GID>
<name>OUT_8</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>560 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-49.5,50.5,-49.5</points>
<connection>
<GID>12</GID>
<name>OUT_9</name></connection>
<connection>
<GID>100</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>254 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-97.5,31,-97.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>272 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-37,23.5,-37</points>
<connection>
<GID>68</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>255 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-96.5,31,-96.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<connection>
<GID>73</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>261 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-87.5,31,-87.5</points>
<connection>
<GID>14</GID>
<name>IN_10</name></connection>
<connection>
<GID>91</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>266 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-86.5,31,-86.5</points>
<connection>
<GID>14</GID>
<name>IN_11</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>262 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-85.5,31,-85.5</points>
<connection>
<GID>14</GID>
<name>IN_12</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>265 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-84.5,31,-84.5</points>
<connection>
<GID>14</GID>
<name>IN_13</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>263 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-83.5,31,-83.5</points>
<connection>
<GID>14</GID>
<name>IN_14</name></connection>
<connection>
<GID>95</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>257 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-94.5,31,-94.5</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<connection>
<GID>77</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>258 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-93.5,31,-93.5</points>
<connection>
<GID>14</GID>
<name>IN_4</name></connection>
<connection>
<GID>85</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>269 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-92.5,31,-92.5</points>
<connection>
<GID>14</GID>
<name>IN_5</name></connection>
<connection>
<GID>86</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>259 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-91.5,31,-91.5</points>
<connection>
<GID>14</GID>
<name>IN_6</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>573 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-83,-5,-80</points>
<connection>
<GID>8</GID>
<name>clear</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-83,-4,-83</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>268 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-90.5,31,-90.5</points>
<connection>
<GID>14</GID>
<name>IN_7</name></connection>
<connection>
<GID>88</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>565 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-42,0,-39</points>
<connection>
<GID>6</GID>
<name>clear</name></connection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>0,-42,1,-42</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>260 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-89.5,31,-89.5</points>
<connection>
<GID>14</GID>
<name>IN_8</name></connection>
<connection>
<GID>89</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>267 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-88.5,31,-88.5</points>
<connection>
<GID>14</GID>
<name>IN_9</name></connection>
<connection>
<GID>90</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>583 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-102.5,37,-99.5</points>
<connection>
<GID>14</GID>
<name>clear</name></connection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-102.5,38,-102.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>496 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-102.5,35,-99.5</points>
<connection>
<GID>14</GID>
<name>clock</name></connection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-102.5,35,-102.5</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>400 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-94.5,41.5,-94.5</points>
<connection>
<GID>14</GID>
<name>OUT_3</name></connection>
<connection>
<GID>55</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>577 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-80.5,36,-77</points>
<connection>
<GID>14</GID>
<name>count_enable</name></connection>
<intersection>-77 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-77,36.5,-77</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>578 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-80.5,37,-80</points>
<connection>
<GID>14</GID>
<name>count_up</name></connection>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>582 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-80.5,35,-79</points>
<connection>
<GID>14</GID>
<name>load</name></connection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-79,35,-79</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>399 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-96.5,41.5,-96.5</points>
<connection>
<GID>14</GID>
<name>OUT_1</name></connection>
<connection>
<GID>55</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>405 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-87.5,41.5,-87.5</points>
<connection>
<GID>14</GID>
<name>OUT_10</name></connection>
<connection>
<GID>55</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>403 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-86.5,41.5,-86.5</points>
<connection>
<GID>14</GID>
<name>OUT_11</name></connection>
<connection>
<GID>55</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>407 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-83.5,41.5,-83.5</points>
<connection>
<GID>14</GID>
<name>OUT_14</name></connection>
<connection>
<GID>55</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>409 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-82.5,41.5,-82.5</points>
<connection>
<GID>14</GID>
<name>OUT_15</name></connection>
<connection>
<GID>55</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>575 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-61,-6,-57.5</points>
<connection>
<GID>8</GID>
<name>count_enable</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-57.5,-5,-57.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>410 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-95.5,41.5,-95.5</points>
<connection>
<GID>14</GID>
<name>OUT_2</name></connection>
<connection>
<GID>55</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>401 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-93.5,41.5,-93.5</points>
<connection>
<GID>14</GID>
<name>OUT_4</name></connection>
<connection>
<GID>55</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>585 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-102,-7.5,-101</points>
<connection>
<GID>16</GID>
<name>load</name></connection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-101,-7.5,-101</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>408 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-92.5,41.5,-92.5</points>
<connection>
<GID>14</GID>
<name>OUT_5</name></connection>
<connection>
<GID>55</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>411 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-91.5,41.5,-91.5</points>
<connection>
<GID>14</GID>
<name>OUT_6</name></connection>
<connection>
<GID>55</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>589 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-144.5,36.5,-141</points>
<connection>
<GID>18</GID>
<name>clear</name></connection>
<intersection>-144.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-144.5,37.5,-144.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>412 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-90.5,41.5,-90.5</points>
<connection>
<GID>14</GID>
<name>OUT_7</name></connection>
<connection>
<GID>55</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>402 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-89.5,41.5,-89.5</points>
<connection>
<GID>14</GID>
<name>OUT_8</name></connection>
<connection>
<GID>55</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>413 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-88.5,41.5,-88.5</points>
<connection>
<GID>14</GID>
<name>OUT_9</name></connection>
<connection>
<GID>55</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>95 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-37,-6,-37</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>179 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-36,-6,-36</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<connection>
<GID>27</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>177 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-27,-6,-27</points>
<connection>
<GID>6</GID>
<name>IN_10</name></connection>
<connection>
<GID>27</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>178 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-26,-6,-26</points>
<connection>
<GID>6</GID>
<name>IN_11</name></connection>
<connection>
<GID>27</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>93 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-35,-6,-35</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<connection>
<GID>27</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>463 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-137,41,-137</points>
<connection>
<GID>18</GID>
<name>OUT_2</name></connection>
<connection>
<GID>59</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>96 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-34,-6,-34</points>
<connection>
<GID>6</GID>
<name>IN_3</name></connection>
<connection>
<GID>27</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>97 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-33,-6,-33</points>
<connection>
<GID>6</GID>
<name>IN_4</name></connection>
<connection>
<GID>27</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>457 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-134,45.5,-134</points>
<connection>
<GID>59</GID>
<name>OUT_5</name></connection>
<connection>
<GID>60</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>98 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-32,-6,-32</points>
<connection>
<GID>6</GID>
<name>IN_5</name></connection>
<connection>
<GID>27</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>176 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-31,-6,-31</points>
<connection>
<GID>6</GID>
<name>IN_6</name></connection>
<connection>
<GID>27</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>453 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-128,45.5,-128</points>
<connection>
<GID>59</GID>
<name>OUT_11</name></connection>
<connection>
<GID>60</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>94 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-30,-6,-30</points>
<connection>
<GID>6</GID>
<name>IN_7</name></connection>
<connection>
<GID>27</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>180 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-29,-6,-29</points>
<connection>
<GID>6</GID>
<name>IN_8</name></connection>
<connection>
<GID>27</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>175 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-28,-6,-28</points>
<connection>
<GID>6</GID>
<name>IN_9</name></connection>
<connection>
<GID>27</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>499 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-42,-2,-39</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3,-42,-2,-42</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>568 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-24,-1,-20.5</points>
<connection>
<GID>6</GID>
<name>count_enable</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1,-20.5,0,-20.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>566 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-24,-2,-22.5</points>
<connection>
<GID>6</GID>
<name>load</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-22.5,-2,-22.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>188 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-37,7,-37</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>182 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-36,7,-36</points>
<connection>
<GID>6</GID>
<name>OUT_1</name></connection>
<connection>
<GID>66</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>191 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-27,7,-27</points>
<connection>
<GID>6</GID>
<name>OUT_10</name></connection>
<connection>
<GID>66</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>192 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-26,7,-26</points>
<connection>
<GID>6</GID>
<name>OUT_11</name></connection>
<connection>
<GID>66</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>190 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-35,7,-35</points>
<connection>
<GID>6</GID>
<name>OUT_2</name></connection>
<connection>
<GID>66</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>189 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-34,7,-34</points>
<connection>
<GID>6</GID>
<name>OUT_3</name></connection>
<connection>
<GID>66</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>181 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-33,7,-33</points>
<connection>
<GID>6</GID>
<name>OUT_4</name></connection>
<connection>
<GID>66</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>183 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-32,7,-32</points>
<connection>
<GID>6</GID>
<name>OUT_5</name></connection>
<connection>
<GID>66</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>184 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-31,7,-31</points>
<connection>
<GID>6</GID>
<name>OUT_6</name></connection>
<connection>
<GID>66</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>185 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-30,7,-30</points>
<connection>
<GID>6</GID>
<name>OUT_7</name></connection>
<connection>
<GID>66</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>187 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-29,7,-29</points>
<connection>
<GID>6</GID>
<name>OUT_8</name></connection>
<connection>
<GID>66</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>186 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-28,7,-28</points>
<connection>
<GID>6</GID>
<name>OUT_9</name></connection>
<connection>
<GID>66</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>125 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-78,-11,-78</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>467 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-138,41,-138</points>
<connection>
<GID>18</GID>
<name>OUT_1</name></connection>
<connection>
<GID>59</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>116 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-77,-11,-77</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>115 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-68,-11,-68</points>
<connection>
<GID>8</GID>
<name>IN_10</name></connection>
<connection>
<GID>34</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>120 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-67,-11,-67</points>
<connection>
<GID>8</GID>
<name>IN_11</name></connection>
<connection>
<GID>34</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>122 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-66,-11,-66</points>
<connection>
<GID>8</GID>
<name>IN_12</name></connection>
<connection>
<GID>34</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>117 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-65,-11,-65</points>
<connection>
<GID>8</GID>
<name>IN_13</name></connection>
<connection>
<GID>34</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>477 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-133,41,-133</points>
<connection>
<GID>18</GID>
<name>OUT_6</name></connection>
<connection>
<GID>59</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>118 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-64,-11,-64</points>
<connection>
<GID>8</GID>
<name>IN_14</name></connection>
<connection>
<GID>34</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>121 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-63,-11,-63</points>
<connection>
<GID>8</GID>
<name>IN_15</name></connection>
<connection>
<GID>34</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>123 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-76,-11,-76</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<connection>
<GID>34</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>112 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-75,-11,-75</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<connection>
<GID>34</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>126 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-74,-11,-74</points>
<connection>
<GID>8</GID>
<name>IN_4</name></connection>
<connection>
<GID>34</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>119 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-73,-11,-73</points>
<connection>
<GID>8</GID>
<name>IN_5</name></connection>
<connection>
<GID>34</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>473 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-130,41,-130</points>
<connection>
<GID>18</GID>
<name>OUT_9</name></connection>
<connection>
<GID>59</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>114 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-72,-11,-72</points>
<connection>
<GID>8</GID>
<name>IN_6</name></connection>
<connection>
<GID>34</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>113 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-71,-11,-71</points>
<connection>
<GID>8</GID>
<name>IN_7</name></connection>
<connection>
<GID>34</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>111 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-70,-11,-70</points>
<connection>
<GID>8</GID>
<name>IN_8</name></connection>
<connection>
<GID>34</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>475 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-134,41,-134</points>
<connection>
<GID>18</GID>
<name>OUT_5</name></connection>
<connection>
<GID>59</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>124 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-69,-11,-69</points>
<connection>
<GID>8</GID>
<name>IN_9</name></connection>
<connection>
<GID>34</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>574 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-61,-5,-60.5</points>
<connection>
<GID>8</GID>
<name>count_up</name></connection>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>369 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-78,-0.5,-78</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>53</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>576 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-61,-7,-59.5</points>
<connection>
<GID>8</GID>
<name>load</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-59.5,-7,-59.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>374 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-77,-0.5,-77</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<connection>
<GID>53</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>377 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-68,-0.5,-68</points>
<connection>
<GID>8</GID>
<name>OUT_10</name></connection>
<connection>
<GID>53</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>379 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-67,-0.5,-67</points>
<connection>
<GID>8</GID>
<name>OUT_11</name></connection>
<connection>
<GID>53</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>588 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-122,34.5,-120.5</points>
<connection>
<GID>18</GID>
<name>load</name></connection>
<intersection>-120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-120.5,34.5,-120.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>381 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-65,-0.5,-65</points>
<connection>
<GID>8</GID>
<name>OUT_13</name></connection>
<connection>
<GID>53</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>371 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-64,-0.5,-64</points>
<connection>
<GID>8</GID>
<name>OUT_14</name></connection>
<connection>
<GID>53</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>382 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-63,-0.5,-63</points>
<connection>
<GID>8</GID>
<name>OUT_15</name></connection>
<connection>
<GID>53</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>375 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-76,-0.5,-76</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<connection>
<GID>53</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>367 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-75,-0.5,-75</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<connection>
<GID>53</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>373 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-74,-0.5,-74</points>
<connection>
<GID>8</GID>
<name>OUT_4</name></connection>
<connection>
<GID>53</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>372 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-73,-0.5,-73</points>
<connection>
<GID>8</GID>
<name>OUT_5</name></connection>
<connection>
<GID>53</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>368 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-72,-0.5,-72</points>
<connection>
<GID>8</GID>
<name>OUT_6</name></connection>
<connection>
<GID>53</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>378 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-71,-0.5,-71</points>
<connection>
<GID>8</GID>
<name>OUT_7</name></connection>
<connection>
<GID>53</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>370 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-70,-0.5,-70</points>
<connection>
<GID>8</GID>
<name>OUT_8</name></connection>
<connection>
<GID>53</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>494 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-144.5,34.5,-141</points>
<connection>
<GID>18</GID>
<name>clock</name></connection>
<intersection>-144.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-144.5,34.5,-144.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>146 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-119,-11.5,-119</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>144 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-118,-11.5,-118</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<connection>
<GID>36</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>147 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-109,-11.5,-109</points>
<connection>
<GID>16</GID>
<name>IN_10</name></connection>
<connection>
<GID>36</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>145 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-108,-11.5,-108</points>
<connection>
<GID>16</GID>
<name>IN_11</name></connection>
<connection>
<GID>36</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>152 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-107,-11.5,-107</points>
<connection>
<GID>16</GID>
<name>IN_12</name></connection>
<connection>
<GID>36</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>153 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-106,-11.5,-106</points>
<connection>
<GID>16</GID>
<name>IN_13</name></connection>
<connection>
<GID>36</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>155 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-105,-11.5,-105</points>
<connection>
<GID>16</GID>
<name>IN_14</name></connection>
<connection>
<GID>36</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>158 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-104,-11.5,-104</points>
<connection>
<GID>16</GID>
<name>IN_15</name></connection>
<connection>
<GID>36</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>150 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-117,-11.5,-117</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<connection>
<GID>36</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>149 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-116,-11.5,-116</points>
<connection>
<GID>16</GID>
<name>IN_3</name></connection>
<connection>
<GID>36</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>148 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-115,-11.5,-115</points>
<connection>
<GID>16</GID>
<name>IN_4</name></connection>
<connection>
<GID>36</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>156 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-114,-11.5,-114</points>
<connection>
<GID>16</GID>
<name>IN_5</name></connection>
<connection>
<GID>36</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>288 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-31,32.5,-31</points>
<connection>
<GID>101</GID>
<name>OUT_6</name></connection>
<connection>
<GID>24</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>143 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-113,-11.5,-113</points>
<connection>
<GID>16</GID>
<name>IN_6</name></connection>
<connection>
<GID>36</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>154 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-112,-11.5,-112</points>
<connection>
<GID>16</GID>
<name>IN_7</name></connection>
<connection>
<GID>36</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>151 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-111,-11.5,-111</points>
<connection>
<GID>16</GID>
<name>IN_8</name></connection>
<connection>
<GID>36</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>157 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-110,-11.5,-110</points>
<connection>
<GID>16</GID>
<name>IN_9</name></connection>
<connection>
<GID>36</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>495 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-124.5,-7.5,-121</points>
<connection>
<GID>16</GID>
<name>clock</name></connection>
<intersection>-124.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,-124.5,-7.5,-124.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>579 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>-5.5,-102,-5.5,-101.5</points>
<connection>
<GID>16</GID>
<name>count_up</name></connection>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>431 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-119,-1,-119</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>439 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-109,-1,-109</points>
<connection>
<GID>16</GID>
<name>OUT_10</name></connection>
<connection>
<GID>57</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>444 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-108,-1,-108</points>
<connection>
<GID>16</GID>
<name>OUT_11</name></connection>
<connection>
<GID>57</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>443 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-107,-1,-107</points>
<connection>
<GID>16</GID>
<name>OUT_12</name></connection>
<connection>
<GID>57</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>445 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-106,-1,-106</points>
<connection>
<GID>16</GID>
<name>OUT_13</name></connection>
<connection>
<GID>57</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>442 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-105,-1,-105</points>
<connection>
<GID>16</GID>
<name>OUT_14</name></connection>
<connection>
<GID>57</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>446 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-104,-1,-104</points>
<connection>
<GID>16</GID>
<name>OUT_15</name></connection>
<connection>
<GID>57</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>433 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-117,-1,-117</points>
<connection>
<GID>16</GID>
<name>OUT_2</name></connection>
<connection>
<GID>57</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>434 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-116,-1,-116</points>
<connection>
<GID>16</GID>
<name>OUT_3</name></connection>
<connection>
<GID>57</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>435 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-115,-1,-115</points>
<connection>
<GID>16</GID>
<name>OUT_4</name></connection>
<connection>
<GID>57</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>440 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-114,-1,-114</points>
<connection>
<GID>16</GID>
<name>OUT_5</name></connection>
<connection>
<GID>57</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>441 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-113,-1,-113</points>
<connection>
<GID>16</GID>
<name>OUT_6</name></connection>
<connection>
<GID>57</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>437 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-111,-1,-111</points>
<connection>
<GID>16</GID>
<name>OUT_8</name></connection>
<connection>
<GID>57</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>438 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-110,-1,-110</points>
<connection>
<GID>16</GID>
<name>OUT_9</name></connection>
<connection>
<GID>57</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>164 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-139,30.5,-139</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>37</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>168 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-138,30.5,-138</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<connection>
<GID>37</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>171 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-129,30.5,-129</points>
<connection>
<GID>18</GID>
<name>IN_10</name></connection>
<connection>
<GID>37</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>172 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-128,30.5,-128</points>
<connection>
<GID>18</GID>
<name>IN_11</name></connection>
<connection>
<GID>37</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>174 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-127,30.5,-127</points>
<connection>
<GID>18</GID>
<name>IN_12</name></connection>
<connection>
<GID>37</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>159 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-126,30.5,-126</points>
<connection>
<GID>18</GID>
<name>IN_13</name></connection>
<connection>
<GID>37</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>162 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-125,30.5,-125</points>
<connection>
<GID>18</GID>
<name>IN_14</name></connection>
<connection>
<GID>37</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>163 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-124,30.5,-124</points>
<connection>
<GID>18</GID>
<name>IN_15</name></connection>
<connection>
<GID>37</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>169 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-137,30.5,-137</points>
<connection>
<GID>18</GID>
<name>IN_2</name></connection>
<connection>
<GID>37</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>165 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-136,30.5,-136</points>
<connection>
<GID>18</GID>
<name>IN_3</name></connection>
<connection>
<GID>37</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>173 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-135,30.5,-135</points>
<connection>
<GID>18</GID>
<name>IN_4</name></connection>
<connection>
<GID>37</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>161 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-134,30.5,-134</points>
<connection>
<GID>18</GID>
<name>IN_5</name></connection>
<connection>
<GID>37</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>167 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-133,30.5,-133</points>
<connection>
<GID>18</GID>
<name>IN_6</name></connection>
<connection>
<GID>37</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>160 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-132,30.5,-132</points>
<connection>
<GID>18</GID>
<name>IN_7</name></connection>
<connection>
<GID>37</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>170 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-131,30.5,-131</points>
<connection>
<GID>18</GID>
<name>IN_8</name></connection>
<connection>
<GID>37</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>166 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-130,30.5,-130</points>
<connection>
<GID>18</GID>
<name>IN_9</name></connection>
<connection>
<GID>37</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>587 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-122,35.5,-118</points>
<connection>
<GID>18</GID>
<name>count_enable</name></connection>
<intersection>-118 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-118,36.5,-118</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>474 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-128,41,-128</points>
<connection>
<GID>18</GID>
<name>OUT_11</name></connection>
<connection>
<GID>59</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>478 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-127,41,-127</points>
<connection>
<GID>18</GID>
<name>OUT_12</name></connection>
<connection>
<GID>59</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>470 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-126,41,-126</points>
<connection>
<GID>18</GID>
<name>OUT_13</name></connection>
<connection>
<GID>59</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>472 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-125,41,-125</points>
<connection>
<GID>18</GID>
<name>OUT_14</name></connection>
<connection>
<GID>59</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>476 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-124,41,-124</points>
<connection>
<GID>18</GID>
<name>OUT_15</name></connection>
<connection>
<GID>59</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>464 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-136,41,-136</points>
<connection>
<GID>18</GID>
<name>OUT_3</name></connection>
<connection>
<GID>59</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>466 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-135,41,-135</points>
<connection>
<GID>18</GID>
<name>OUT_4</name></connection>
<connection>
<GID>59</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>468 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-132,41,-132</points>
<connection>
<GID>18</GID>
<name>OUT_7</name></connection>
<connection>
<GID>59</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>294 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-37,32.5,-37</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>293 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-36,32.5,-36</points>
<connection>
<GID>101</GID>
<name>OUT_1</name></connection>
<connection>
<GID>24</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>282 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32,-27,32.5,-27</points>
<connection>
<GID>102</GID>
<name>OUT_2</name></connection>
<connection>
<GID>24</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>292 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-35,32.5,-35</points>
<connection>
<GID>101</GID>
<name>OUT_2</name></connection>
<connection>
<GID>24</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>291 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-34,32.5,-34</points>
<connection>
<GID>101</GID>
<name>OUT_3</name></connection>
<connection>
<GID>24</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>290 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-33,32.5,-33</points>
<connection>
<GID>101</GID>
<name>OUT_4</name></connection>
<connection>
<GID>24</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>289 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-32,32.5,-32</points>
<connection>
<GID>101</GID>
<name>OUT_5</name></connection>
<connection>
<GID>24</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>287 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-30,32.5,-30</points>
<connection>
<GID>101</GID>
<name>OUT_7</name></connection>
<connection>
<GID>24</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>279 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32,-29,32.5,-29</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>280 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32,-28,32.5,-28</points>
<connection>
<GID>102</GID>
<name>OUT_1</name></connection>
<connection>
<GID>24</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-7,23,-3</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>-7 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-24.5,-163,-24.5,-7</points>
<intersection>-163 8</intersection>
<intersection>-144 16</intersection>
<intersection>-131.5 34</intersection>
<intersection>-111.5 37</intersection>
<intersection>-70.5 48</intersection>
<intersection>-51 6</intersection>
<intersection>-29.5 55</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24.5,-7,23,-7</points>
<intersection>-24.5 1</intersection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-24.5,-51,22.5,-51</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-24.5,-163,67.5,-163</points>
<intersection>-24.5 1</intersection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-24.5,-144,-13.5,-144</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>67.5,-163,67.5,-29.5</points>
<intersection>-163 8</intersection>
<intersection>-131.5 39</intersection>
<intersection>-111.5 38</intersection>
<intersection>-90 44</intersection>
<intersection>-70.5 50</intersection>
<intersection>-51 49</intersection>
<intersection>-29.5 52</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>-24.5,-131.5,26,-131.5</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-24.5,-111.5,-16,-111.5</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>7.5,-111.5,67.5,-111.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>49.5,-131.5,67.5,-131.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>50,-90,67.5,-90</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-24.5,-70.5,-15.5,-70.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>63.5,-51,67.5,-51</points>
<connection>
<GID>137</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>8,-70.5,67.5,-70.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>36.5,-29.5,67.5,-29.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>-24.5,-29.5,-17.5,-29.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>391 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-82.5,46,-82.5</points>
<connection>
<GID>55</GID>
<name>OUT_15</name></connection>
<connection>
<GID>56</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>385 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-90.5,46,-90.5</points>
<connection>
<GID>55</GID>
<name>OUT_7</name></connection>
<connection>
<GID>56</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>389 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-86.5,46,-86.5</points>
<connection>
<GID>55</GID>
<name>OUT_11</name></connection>
<connection>
<GID>56</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>388 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-83.5,46,-83.5</points>
<connection>
<GID>55</GID>
<name>OUT_14</name></connection>
<connection>
<GID>56</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>693 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-46,52.5,-40</points>
<connection>
<GID>100</GID>
<name>ENABLE_0</name></connection>
<intersection>-46 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-40,53.5,-40</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-46,52.5,-46</points>
<intersection>48 8</intersection>
<intersection>52.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>48,-50,48,-46</points>
<connection>
<GID>99</GID>
<name>ENABLE_0</name></connection>
<intersection>-46 2</intersection></vsegment></shape></wire>
<wire>
<ID>661 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-58.5,59.5,-58.5</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<connection>
<GID>137</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>662 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-57.5,59.5,-57.5</points>
<connection>
<GID>99</GID>
<name>OUT_1</name></connection>
<connection>
<GID>137</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>663 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-56.5,59.5,-56.5</points>
<connection>
<GID>99</GID>
<name>OUT_2</name></connection>
<connection>
<GID>137</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>664 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-55.5,59.5,-55.5</points>
<connection>
<GID>99</GID>
<name>OUT_3</name></connection>
<connection>
<GID>137</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>665 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-54.5,59.5,-54.5</points>
<connection>
<GID>99</GID>
<name>OUT_4</name></connection>
<connection>
<GID>137</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>666 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-53.5,59.5,-53.5</points>
<connection>
<GID>99</GID>
<name>OUT_5</name></connection>
<connection>
<GID>137</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>667 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-52.5,59.5,-52.5</points>
<connection>
<GID>99</GID>
<name>OUT_6</name></connection>
<connection>
<GID>137</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>668 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-51.5,59.5,-51.5</points>
<connection>
<GID>99</GID>
<name>OUT_7</name></connection>
<connection>
<GID>137</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>657 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-50.5,59.5,-50.5</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<connection>
<GID>137</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>658 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-49.5,59.5,-49.5</points>
<connection>
<GID>100</GID>
<name>OUT_1</name></connection>
<connection>
<GID>137</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>660 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-48.5,59.5,-48.5</points>
<connection>
<GID>100</GID>
<name>OUT_2</name></connection>
<connection>
<GID>137</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>659 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-47.5,59.5,-47.5</points>
<connection>
<GID>100</GID>
<name>OUT_3</name></connection>
<connection>
<GID>137</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>694 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-61.5,1.5,-59.5</points>
<connection>
<GID>53</GID>
<name>ENABLE_0</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1.5,-59.5,6,-59.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>365 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-78,4,-78</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<connection>
<GID>54</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>366 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-77,4,-77</points>
<connection>
<GID>53</GID>
<name>OUT_1</name></connection>
<connection>
<GID>54</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>352 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-68,4,-68</points>
<connection>
<GID>53</GID>
<name>OUT_10</name></connection>
<connection>
<GID>54</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>357 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-67,4,-67</points>
<connection>
<GID>53</GID>
<name>OUT_11</name></connection>
<connection>
<GID>54</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>351 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-66,4,-66</points>
<connection>
<GID>53</GID>
<name>OUT_12</name></connection>
<connection>
<GID>54</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-13,3.5,14.5</points>
<intersection>-13 1</intersection>
<intersection>14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-13,15.5,-13</points>
<intersection>3.5 0</intersection>
<intersection>15.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,14.5,8.5,14.5</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>3.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15.5,-29.5,15.5,-13</points>
<intersection>-29.5 4</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>11,-29.5,18.5,-29.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>15.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>358 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-65,4,-65</points>
<connection>
<GID>53</GID>
<name>OUT_13</name></connection>
<connection>
<GID>54</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>359 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-63,4,-63</points>
<connection>
<GID>53</GID>
<name>OUT_15</name></connection>
<connection>
<GID>54</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>362 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-76,4,-76</points>
<connection>
<GID>53</GID>
<name>OUT_2</name></connection>
<connection>
<GID>54</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>363 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-75,4,-75</points>
<connection>
<GID>53</GID>
<name>OUT_3</name></connection>
<connection>
<GID>54</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>360 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-74,4,-74</points>
<connection>
<GID>53</GID>
<name>OUT_4</name></connection>
<connection>
<GID>54</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>696 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-102.5,1,-100.5</points>
<connection>
<GID>57</GID>
<name>ENABLE_0</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-100.5,5,-100.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>361 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-73,4,-73</points>
<connection>
<GID>53</GID>
<name>OUT_5</name></connection>
<connection>
<GID>54</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>353 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-71,4,-71</points>
<connection>
<GID>53</GID>
<name>OUT_7</name></connection>
<connection>
<GID>54</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>355 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-69,4,-69</points>
<connection>
<GID>53</GID>
<name>OUT_9</name></connection>
<connection>
<GID>54</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>695 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-81,43.5,-79</points>
<connection>
<GID>55</GID>
<name>ENABLE_0</name></connection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-79,49.5,-79</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>397 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-97.5,46,-97.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<connection>
<GID>56</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>398 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-96.5,46,-96.5</points>
<connection>
<GID>55</GID>
<name>OUT_1</name></connection>
<connection>
<GID>56</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>384 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-87.5,46,-87.5</points>
<connection>
<GID>55</GID>
<name>OUT_10</name></connection>
<connection>
<GID>56</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>383 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-85.5,46,-85.5</points>
<connection>
<GID>55</GID>
<name>OUT_12</name></connection>
<connection>
<GID>56</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>390 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-84.5,46,-84.5</points>
<connection>
<GID>55</GID>
<name>OUT_13</name></connection>
<connection>
<GID>56</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>395 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-94.5,46,-94.5</points>
<connection>
<GID>55</GID>
<name>OUT_3</name></connection>
<connection>
<GID>56</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>697 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-122.5,43,-119.5</points>
<connection>
<GID>59</GID>
<name>ENABLE_0</name></connection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>43,-119.5,46,-119.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>392 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-93.5,46,-93.5</points>
<connection>
<GID>55</GID>
<name>OUT_4</name></connection>
<connection>
<GID>56</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>393 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-92.5,46,-92.5</points>
<connection>
<GID>55</GID>
<name>OUT_5</name></connection>
<connection>
<GID>56</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>396 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-91.5,46,-91.5</points>
<connection>
<GID>55</GID>
<name>OUT_6</name></connection>
<connection>
<GID>56</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>387 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-88.5,46,-88.5</points>
<connection>
<GID>55</GID>
<name>OUT_9</name></connection>
<connection>
<GID>56</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>429 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-119,3.5,-119</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<connection>
<GID>58</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>430 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-118,3.5,-118</points>
<connection>
<GID>57</GID>
<name>OUT_1</name></connection>
<connection>
<GID>58</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>416 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-109,3.5,-109</points>
<connection>
<GID>57</GID>
<name>OUT_10</name></connection>
<connection>
<GID>58</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>421 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-108,3.5,-108</points>
<connection>
<GID>57</GID>
<name>OUT_11</name></connection>
<connection>
<GID>58</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>415 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-107,3.5,-107</points>
<connection>
<GID>57</GID>
<name>OUT_12</name></connection>
<connection>
<GID>58</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>420 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-105,3.5,-105</points>
<connection>
<GID>57</GID>
<name>OUT_14</name></connection>
<connection>
<GID>58</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>423 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-104,3.5,-104</points>
<connection>
<GID>57</GID>
<name>OUT_15</name></connection>
<connection>
<GID>58</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>426 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-117,3.5,-117</points>
<connection>
<GID>57</GID>
<name>OUT_2</name></connection>
<connection>
<GID>58</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>427 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-116,3.5,-116</points>
<connection>
<GID>57</GID>
<name>OUT_3</name></connection>
<connection>
<GID>58</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>424 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-115,3.5,-115</points>
<connection>
<GID>57</GID>
<name>OUT_4</name></connection>
<connection>
<GID>58</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>425 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-114,3.5,-114</points>
<connection>
<GID>57</GID>
<name>OUT_5</name></connection>
<connection>
<GID>58</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>428 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-113,3.5,-113</points>
<connection>
<GID>57</GID>
<name>OUT_6</name></connection>
<connection>
<GID>58</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>418 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-111,3.5,-111</points>
<connection>
<GID>57</GID>
<name>OUT_8</name></connection>
<connection>
<GID>58</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>419 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-110,3.5,-110</points>
<connection>
<GID>57</GID>
<name>OUT_9</name></connection>
<connection>
<GID>58</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>417 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-112,3.5,-112</points>
<connection>
<GID>57</GID>
<name>OUT_7</name></connection>
<connection>
<GID>58</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>448 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-129,45.5,-129</points>
<connection>
<GID>59</GID>
<name>OUT_10</name></connection>
<connection>
<GID>60</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>447 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-127,45.5,-127</points>
<connection>
<GID>59</GID>
<name>OUT_12</name></connection>
<connection>
<GID>60</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>454 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-126,45.5,-126</points>
<connection>
<GID>59</GID>
<name>OUT_13</name></connection>
<connection>
<GID>60</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>452 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-125,45.5,-125</points>
<connection>
<GID>59</GID>
<name>OUT_14</name></connection>
<connection>
<GID>60</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>455 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-124,45.5,-124</points>
<connection>
<GID>59</GID>
<name>OUT_15</name></connection>
<connection>
<GID>60</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>458 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-137,45.5,-137</points>
<connection>
<GID>59</GID>
<name>OUT_2</name></connection>
<connection>
<GID>60</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>456 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-135,45.5,-135</points>
<connection>
<GID>59</GID>
<name>OUT_4</name></connection>
<connection>
<GID>60</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>460 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-133,45.5,-133</points>
<connection>
<GID>59</GID>
<name>OUT_6</name></connection>
<connection>
<GID>60</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>449 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-132,45.5,-132</points>
<connection>
<GID>59</GID>
<name>OUT_7</name></connection>
<connection>
<GID>60</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>276 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-36,23.5,-36</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<connection>
<GID>101</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>285 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-27,28,-27</points>
<connection>
<GID>68</GID>
<name>IN_10</name></connection>
<connection>
<GID>102</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>286 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-26,28,-26</points>
<connection>
<GID>68</GID>
<name>IN_11</name></connection>
<connection>
<GID>102</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>273 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-35,23.5,-35</points>
<connection>
<GID>68</GID>
<name>IN_2</name></connection>
<connection>
<GID>101</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>275 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-34,23.5,-34</points>
<connection>
<GID>68</GID>
<name>IN_3</name></connection>
<connection>
<GID>101</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>271 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-32,23.5,-32</points>
<connection>
<GID>68</GID>
<name>IN_5</name></connection>
<connection>
<GID>101</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>274 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-31,23.5,-31</points>
<connection>
<GID>68</GID>
<name>IN_6</name></connection>
<connection>
<GID>101</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>278 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-30,23.5,-30</points>
<connection>
<GID>68</GID>
<name>IN_7</name></connection>
<connection>
<GID>101</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>283 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-29,28,-29</points>
<connection>
<GID>68</GID>
<name>IN_8</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>284 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-28,28,-28</points>
<connection>
<GID>68</GID>
<name>IN_9</name></connection>
<connection>
<GID>102</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>295 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-24.5,30,-18</points>
<connection>
<GID>102</GID>
<name>ENABLE_0</name></connection>
<intersection>-24.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-18,31,-18</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-24.5,30,-24.5</points>
<intersection>25.5 3</intersection>
<intersection>30 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25.5,-28.5,25.5,-24.5</points>
<connection>
<GID>101</GID>
<name>ENABLE_0</name></connection>
<intersection>-24.5 2</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-176.453,80.375,312.403,-166.25</PageViewport>
<gate>
<ID>310</ID>
<type>AA_AND2</type>
<position>96,-20</position>
<input>
<ID>IN_0</ID>511 </input>
<input>
<ID>IN_1</ID>510 </input>
<output>
<ID>OUT</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>DA_FROM</type>
<position>13,70.5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND2</type>
<position>-50,-40</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>AE_FULLADDER_4BIT</type>
<position>21.5,17</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>132 </input>
<input>
<ID>IN_2</ID>130 </input>
<input>
<ID>IN_3</ID>131 </input>
<input>
<ID>IN_B_0</ID>226 </input>
<input>
<ID>IN_B_1</ID>225 </input>
<input>
<ID>IN_B_2</ID>224 </input>
<input>
<ID>IN_B_3</ID>223 </input>
<output>
<ID>OUT_0</ID>243 </output>
<output>
<ID>OUT_1</ID>241 </output>
<output>
<ID>OUT_2</ID>242 </output>
<output>
<ID>OUT_3</ID>244 </output>
<input>
<ID>carry_in</ID>77 </input>
<output>
<ID>carry_out</ID>81 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_AND2</type>
<position>-50,-15</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>-70,-39</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>-50,-10</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_AND2</type>
<position>-64.5,-11</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>AE_FULLADDER_4BIT</type>
<position>21.5,53</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>90 </input>
<input>
<ID>IN_2</ID>88 </input>
<input>
<ID>IN_3</ID>89 </input>
<input>
<ID>IN_B_0</ID>140 </input>
<input>
<ID>IN_B_1</ID>139 </input>
<input>
<ID>IN_B_2</ID>138 </input>
<input>
<ID>IN_B_3</ID>137 </input>
<output>
<ID>OUT_0</ID>233 </output>
<output>
<ID>OUT_1</ID>234 </output>
<output>
<ID>OUT_2</ID>235 </output>
<output>
<ID>OUT_3</ID>236 </output>
<input>
<ID>carry_in</ID>78 </input>
<output>
<ID>carry_out</ID>79 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>509</ID>
<type>AA_AND2</type>
<position>23,-123</position>
<input>
<ID>IN_0</ID>755 </input>
<input>
<ID>IN_1</ID>756 </input>
<output>
<ID>OUT</ID>739 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>-50,-20</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>DA_FROM</type>
<position>13,66.5</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>-70,-7</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>151</ID>
<type>AE_FULLADDER_4BIT</type>
<position>21.5,71</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>84 </input>
<input>
<ID>IN_2</ID>85 </input>
<input>
<ID>IN_3</ID>86 </input>
<input>
<ID>IN_B_0</ID>133 </input>
<input>
<ID>IN_B_1</ID>134 </input>
<input>
<ID>IN_B_2</ID>135 </input>
<input>
<ID>IN_B_3</ID>136 </input>
<output>
<ID>OUT_0</ID>231 </output>
<output>
<ID>OUT_1</ID>228 </output>
<output>
<ID>OUT_2</ID>230 </output>
<output>
<ID>OUT_3</ID>232 </output>
<input>
<ID>carry_in</ID>82 </input>
<output>
<ID>carry_out</ID>78 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND2</type>
<position>-50,-25</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>154</ID>
<type>DE_TO</type>
<position>33.5,5</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cout</lparam></gate>
<gate>
<ID>385</ID>
<type>DA_FROM</type>
<position>149,-57</position>
<input>
<ID>IN_0</ID>708 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add7</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND2</type>
<position>-50,-30</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>FF_GND</type>
<position>26.5,78</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>507</ID>
<type>DA_FROM</type>
<position>-70,-134</position>
<input>
<ID>IN_0</ID>811 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND2</type>
<position>-50,-35</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>13,48.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>-70,-10</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>397</ID>
<type>AA_AND2</type>
<position>23,-66</position>
<input>
<ID>IN_0</ID>631 </input>
<input>
<ID>IN_1</ID>632 </input>
<output>
<ID>OUT</ID>625 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>-70,-12</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>-70,-14</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>173</ID>
<type>DA_FROM</type>
<position>13,28.5</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_OR8</type>
<position>-21.5,-25.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>41 </input>
<input>
<ID>IN_4</ID>38 </input>
<input>
<ID>IN_5</ID>38 </input>
<input>
<ID>IN_6</ID>39 </input>
<input>
<ID>IN_7</ID>40 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>174</ID>
<type>DA_FROM</type>
<position>13,16.5</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>469</ID>
<type>AA_AND2</type>
<position>-50,-108</position>
<input>
<ID>IN_0</ID>723 </input>
<input>
<ID>IN_1</ID>724 </input>
<output>
<ID>OUT</ID>717 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>DD_KEYPAD_HEX</type>
<position>56.5,49.5</position>
<output>
<ID>OUT_0</ID>63 </output>
<output>
<ID>OUT_1</ID>64 </output>
<output>
<ID>OUT_2</ID>65 </output>
<output>
<ID>OUT_3</ID>66 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>405</ID>
<type>DA_FROM</type>
<position>3,-62</position>
<input>
<ID>IN_0</ID>629 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>46</ID>
<type>DA_FROM</type>
<position>-70,-19</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>13,14.5</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>47</ID>
<type>DA_FROM</type>
<position>-70,-21</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>13,12.5</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>415</ID>
<type>DA_FROM</type>
<position>3,-57</position>
<input>
<ID>IN_0</ID>641 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add5</lparam></gate>
<gate>
<ID>48</ID>
<type>DA_FROM</type>
<position>-70,-24</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>13,10.5</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>49</ID>
<type>DA_FROM</type>
<position>-70,-26</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp0</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>13,79</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>409</ID>
<type>DA_FROM</type>
<position>3,-72</position>
<input>
<ID>IN_0</ID>634 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>-70,-29</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>179</ID>
<type>DA_FROM</type>
<position>13,75</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>51</ID>
<type>DA_FROM</type>
<position>-70,-31</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_SMALL_INVERTER</type>
<position>-61.5,-31</position>
<input>
<ID>IN_0</ID>51 </input>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>-70,-34</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>129</ID>
<type>DA_FROM</type>
<position>65,30</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>-70,-36</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>70</ID>
<type>DA_FROM</type>
<position>-70,-41</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>471</ID>
<type>AA_AND2</type>
<position>-50,-113</position>
<input>
<ID>IN_0</ID>725 </input>
<input>
<ID>IN_1</ID>727 </input>
<output>
<ID>OUT</ID>716 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AE_REGISTER8</type>
<position>69,43</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>60 </input>
<input>
<ID>IN_4</ID>63 </input>
<input>
<ID>IN_5</ID>64 </input>
<input>
<ID>IN_6</ID>65 </input>
<input>
<ID>IN_7</ID>66 </input>
<output>
<ID>OUT_0</ID>75 </output>
<output>
<ID>OUT_1</ID>74 </output>
<output>
<ID>OUT_2</ID>73 </output>
<output>
<ID>OUT_3</ID>72 </output>
<output>
<ID>OUT_4</ID>71 </output>
<output>
<ID>OUT_5</ID>70 </output>
<output>
<ID>OUT_6</ID>69 </output>
<output>
<ID>OUT_7</ID>68 </output>
<input>
<ID>clock</ID>67 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>123</ID>
<type>DD_KEYPAD_HEX</type>
<position>56.5,37.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<output>
<ID>OUT_1</ID>58 </output>
<output>
<ID>OUT_2</ID>59 </output>
<output>
<ID>OUT_3</ID>60 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>135</ID>
<type>DE_TO</type>
<position>79,47</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp7</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_TO</type>
<position>86.5,46</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp6</lparam></gate>
<gate>
<ID>139</ID>
<type>DE_TO</type>
<position>79,45</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp5</lparam></gate>
<gate>
<ID>140</ID>
<type>DE_TO</type>
<position>86.5,44</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp4</lparam></gate>
<gate>
<ID>141</ID>
<type>DE_TO</type>
<position>79,43</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp3</lparam></gate>
<gate>
<ID>142</ID>
<type>DE_TO</type>
<position>86.5,42</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp2</lparam></gate>
<gate>
<ID>143</ID>
<type>DE_TO</type>
<position>79,41</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp1</lparam></gate>
<gate>
<ID>144</ID>
<type>DE_TO</type>
<position>86.5,40</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp0</lparam></gate>
<gate>
<ID>145</ID>
<type>DE_TO</type>
<position>-13.5,-25.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0in</lparam></gate>
<gate>
<ID>148</ID>
<type>AE_FULLADDER_4BIT</type>
<position>21.5,35</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>92 </input>
<input>
<ID>IN_2</ID>127 </input>
<input>
<ID>IN_3</ID>128 </input>
<input>
<ID>IN_B_0</ID>222 </input>
<input>
<ID>IN_B_1</ID>221 </input>
<input>
<ID>IN_B_2</ID>142 </input>
<input>
<ID>IN_B_3</ID>141 </input>
<output>
<ID>OUT_0</ID>237 </output>
<output>
<ID>OUT_1</ID>238 </output>
<output>
<ID>OUT_2</ID>239 </output>
<output>
<ID>OUT_3</ID>240 </output>
<input>
<ID>carry_in</ID>79 </input>
<output>
<ID>carry_out</ID>77 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>152</ID>
<type>AE_SMALL_INVERTER</type>
<position>27,3</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>306</ID>
<type>AA_AND2</type>
<position>96,-15</position>
<input>
<ID>IN_0</ID>502 </input>
<input>
<ID>IN_1</ID>522 </input>
<output>
<ID>OUT</ID>508 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>DE_TO</type>
<position>33.5,3</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /cout</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>13,68.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>13,64.5</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>314</ID>
<type>AA_AND2</type>
<position>96,-35</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>518 </input>
<output>
<ID>OUT</ID>504 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>DA_FROM</type>
<position>13,52.5</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>162</ID>
<type>DA_FROM</type>
<position>13,50.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>169</ID>
<type>DA_FROM</type>
<position>13,46.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>170</ID>
<type>DA_FROM</type>
<position>13,34.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>171</ID>
<type>DA_FROM</type>
<position>13,32.5</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>13,30.5</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>186</ID>
<type>DA_FROM</type>
<position>13,77</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>187</ID>
<type>DA_FROM</type>
<position>13,73</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>194</ID>
<type>DA_FROM</type>
<position>13,61</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>533</ID>
<type>DA_FROM</type>
<position>3,-119</position>
<input>
<ID>IN_0</ID>754 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>356</ID>
<type>DA_FROM</type>
<position>149,-16</position>
<input>
<ID>IN_0</ID>547 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add3</lparam></gate>
<gate>
<ID>195</ID>
<type>DA_FROM</type>
<position>13,57</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>526</ID>
<type>DA_FROM</type>
<position>3,-104</position>
<input>
<ID>IN_0</ID>746 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>196</ID>
<type>DA_FROM</type>
<position>13,59</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>350</ID>
<type>DA_FROM</type>
<position>149,-31</position>
<input>
<ID>IN_0</ID>540 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>197</ID>
<type>DA_FROM</type>
<position>13,55</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>198</ID>
<type>DA_FROM</type>
<position>13,43</position>
<input>
<ID>IN_0</ID>222 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>521</ID>
<type>DA_FROM</type>
<position>3,-93</position>
<input>
<ID>IN_0</ID>736 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>344</ID>
<type>DE_OR8</type>
<position>197.5,-25.5</position>
<input>
<ID>IN_0</ID>534 </input>
<input>
<ID>IN_1</ID>533 </input>
<input>
<ID>IN_2</ID>532 </input>
<input>
<ID>IN_3</ID>531 </input>
<input>
<ID>IN_4</ID>528 </input>
<input>
<ID>IN_5</ID>528 </input>
<input>
<ID>IN_6</ID>529 </input>
<input>
<ID>IN_7</ID>530 </input>
<output>
<ID>OUT</ID>546 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>199</ID>
<type>DA_FROM</type>
<position>13,39</position>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>530</ID>
<type>DA_FROM</type>
<position>3,-114</position>
<input>
<ID>IN_0</ID>751 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>200</ID>
<type>DA_FROM</type>
<position>13,41</position>
<input>
<ID>IN_0</ID>221 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>354</ID>
<type>DA_FROM</type>
<position>149,-41</position>
<input>
<ID>IN_0</ID>545 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>201</ID>
<type>DA_FROM</type>
<position>13,37</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>202</ID>
<type>DA_FROM</type>
<position>13,25</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>541</ID>
<type>DA_FROM</type>
<position>76,-90</position>
<input>
<ID>IN_0</ID>760 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>364</ID>
<type>DA_FROM</type>
<position>-70,-48</position>
<input>
<ID>IN_0</ID>549 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>203</ID>
<type>DA_FROM</type>
<position>13,21</position>
<input>
<ID>IN_0</ID>224 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>534</ID>
<type>DA_FROM</type>
<position>3,-124</position>
<input>
<ID>IN_0</ID>756 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>204</ID>
<type>DA_FROM</type>
<position>13,23</position>
<input>
<ID>IN_0</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>358</ID>
<type>AA_AND2</type>
<position>-50,-81</position>
<input>
<ID>IN_0</ID>605 </input>
<input>
<ID>IN_1</ID>606 </input>
<output>
<ID>OUT</ID>584 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>DA_FROM</type>
<position>13,19</position>
<input>
<ID>IN_0</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>210</ID>
<type>DA_FROM</type>
<position>-70,-16</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add0</lparam></gate>
<gate>
<ID>549</ID>
<type>DA_FROM</type>
<position>76,-104</position>
<input>
<ID>IN_0</ID>771 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>372</ID>
<type>DA_FROM</type>
<position>-70,-60</position>
<input>
<ID>IN_0</ID>597 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>211</ID>
<type>DE_TO</type>
<position>30,74</position>
<input>
<ID>IN_0</ID>231 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add0</lparam></gate>
<gate>
<ID>542</ID>
<type>AA_AND2</type>
<position>96,-108</position>
<input>
<ID>IN_0</ID>773 </input>
<input>
<ID>IN_1</ID>774 </input>
<output>
<ID>OUT</ID>767 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>DE_TO</type>
<position>30,72</position>
<input>
<ID>IN_0</ID>228 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add1</lparam></gate>
<gate>
<ID>366</ID>
<type>AA_AND2</type>
<position>-50,-71</position>
<input>
<ID>IN_0</ID>600 </input>
<input>
<ID>IN_1</ID>602 </input>
<output>
<ID>OUT</ID>590 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>DE_TO</type>
<position>30,70</position>
<input>
<ID>IN_0</ID>230 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add2</lparam></gate>
<gate>
<ID>214</ID>
<type>DE_TO</type>
<position>30,68</position>
<input>
<ID>IN_0</ID>232 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add3</lparam></gate>
<gate>
<ID>537</ID>
<type>AA_AND2</type>
<position>96,-123</position>
<input>
<ID>IN_0</ID>780 </input>
<input>
<ID>IN_1</ID>781 </input>
<output>
<ID>OUT</ID>764 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>360</ID>
<type>DA_FROM</type>
<position>-70,-80</position>
<input>
<ID>IN_0</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>215</ID>
<type>DE_TO</type>
<position>30,56</position>
<input>
<ID>IN_0</ID>233 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add4</lparam></gate>
<gate>
<ID>546</ID>
<type>DA_FROM</type>
<position>76,-97</position>
<input>
<ID>IN_0</ID>763 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>216</ID>
<type>DE_TO</type>
<position>30,54</position>
<input>
<ID>IN_0</ID>234 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add5</lparam></gate>
<gate>
<ID>370</ID>
<type>DA_FROM</type>
<position>-70,-55</position>
<input>
<ID>IN_0</ID>580 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>217</ID>
<type>DE_TO</type>
<position>30,52</position>
<input>
<ID>IN_0</ID>235 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add6</lparam></gate>
<gate>
<ID>218</ID>
<type>DE_TO</type>
<position>30,50</position>
<input>
<ID>IN_0</ID>236 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add7</lparam></gate>
<gate>
<ID>557</ID>
<type>DA_FROM</type>
<position>76,-124</position>
<input>
<ID>IN_0</ID>781 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>380</ID>
<type>DA_FROM</type>
<position>-70,-77</position>
<input>
<ID>IN_0</ID>604 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>219</ID>
<type>DE_TO</type>
<position>30,38</position>
<input>
<ID>IN_0</ID>237 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add8</lparam></gate>
<gate>
<ID>550</ID>
<type>DA_FROM</type>
<position>76,-107</position>
<input>
<ID>IN_0</ID>773 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>220</ID>
<type>DE_TO</type>
<position>30,36</position>
<input>
<ID>IN_0</ID>238 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add9</lparam></gate>
<gate>
<ID>374</ID>
<type>DA_FROM</type>
<position>-70,-65</position>
<input>
<ID>IN_0</ID>598 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>221</ID>
<type>DE_TO</type>
<position>30,34</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add10</lparam></gate>
<gate>
<ID>222</ID>
<type>DE_TO</type>
<position>30,32</position>
<input>
<ID>IN_0</ID>240 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add11</lparam></gate>
<gate>
<ID>545</ID>
<type>DA_FROM</type>
<position>76,-95</position>
<input>
<ID>IN_0</ID>762 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>368</ID>
<type>DA_FROM</type>
<position>-70,-51</position>
<input>
<ID>IN_0</ID>550 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>223</ID>
<type>DE_TO</type>
<position>30,20</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add12</lparam></gate>
<gate>
<ID>554</ID>
<type>AE_SMALL_INVERTER</type>
<position>84.5,-114</position>
<input>
<ID>IN_0</ID>776 </input>
<output>
<ID>OUT_0</ID>777 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>224</ID>
<type>DE_TO</type>
<position>30,18</position>
<input>
<ID>IN_0</ID>241 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add13</lparam></gate>
<gate>
<ID>378</ID>
<type>AE_SMALL_INVERTER</type>
<position>-61.5,-72</position>
<input>
<ID>IN_0</ID>601 </input>
<output>
<ID>OUT_0</ID>602 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>225</ID>
<type>DE_TO</type>
<position>30,16</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add14</lparam></gate>
<gate>
<ID>226</ID>
<type>DE_TO</type>
<position>30,14</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add15</lparam></gate>
<gate>
<ID>565</ID>
<type>AA_AND2</type>
<position>169,-103</position>
<input>
<ID>IN_0</ID>797 </input>
<input>
<ID>IN_1</ID>796 </input>
<output>
<ID>OUT</ID>793 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_AND2</type>
<position>23,-40</position>
<input>
<ID>IN_0</ID>307 </input>
<input>
<ID>IN_1</ID>308 </input>
<output>
<ID>OUT</ID>250 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>558</ID>
<type>DE_TO</type>
<position>132.5,-108.5</position>
<input>
<ID>IN_0</ID>782 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10in</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_AND2</type>
<position>23,-15</position>
<input>
<ID>IN_0</ID>249 </input>
<input>
<ID>IN_1</ID>310 </input>
<output>
<ID>OUT</ID>296 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>382</ID>
<type>DE_TO</type>
<position>-13.5,-66.5</position>
<input>
<ID>IN_0</ID>607 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4in</lparam></gate>
<gate>
<ID>229</ID>
<type>DA_FROM</type>
<position>3,-39</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_AND2</type>
<position>23,-10</position>
<input>
<ID>IN_0</ID>246 </input>
<input>
<ID>IN_1</ID>245 </input>
<output>
<ID>OUT</ID>297 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>553</ID>
<type>DA_FROM</type>
<position>76,-114</position>
<input>
<ID>IN_0</ID>776 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>376</ID>
<type>DA_FROM</type>
<position>-70,-70</position>
<input>
<ID>IN_0</ID>600 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>231</ID>
<type>AA_AND2</type>
<position>8.5,-11</position>
<input>
<ID>IN_0</ID>247 </input>
<input>
<ID>IN_1</ID>248 </input>
<output>
<ID>OUT</ID>245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>562</ID>
<type>DA_FROM</type>
<position>149,-122</position>
<input>
<ID>IN_0</ID>805 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_AND2</type>
<position>23,-20</position>
<input>
<ID>IN_0</ID>299 </input>
<input>
<ID>IN_1</ID>298 </input>
<output>
<ID>OUT</ID>270 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>233</ID>
<type>DA_FROM</type>
<position>3,-7</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>234</ID>
<type>AA_AND2</type>
<position>23,-25</position>
<input>
<ID>IN_0</ID>300 </input>
<input>
<ID>IN_1</ID>301 </input>
<output>
<ID>OUT</ID>253 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>573</ID>
<type>DA_FROM</type>
<position>149,-102</position>
<input>
<ID>IN_0</ID>797 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>235</ID>
<type>AA_AND2</type>
<position>23,-30</position>
<input>
<ID>IN_0</ID>302 </input>
<input>
<ID>IN_1</ID>304 </input>
<output>
<ID>OUT</ID>252 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>566</ID>
<type>DA_FROM</type>
<position>149,-90</position>
<input>
<ID>IN_0</ID>785 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>23,-35</position>
<input>
<ID>IN_0</ID>305 </input>
<input>
<ID>IN_1</ID>306 </input>
<output>
<ID>OUT</ID>251 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>DA_FROM</type>
<position>3,-10</position>
<input>
<ID>IN_0</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>238</ID>
<type>DA_FROM</type>
<position>3,-12</position>
<input>
<ID>IN_0</ID>248 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>561</ID>
<type>AA_AND2</type>
<position>169,-98</position>
<input>
<ID>IN_0</ID>788 </input>
<input>
<ID>IN_1</ID>808 </input>
<output>
<ID>OUT</ID>794 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>DA_FROM</type>
<position>3,-14</position>
<input>
<ID>IN_0</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>570</ID>
<type>DA_FROM</type>
<position>149,-93</position>
<input>
<ID>IN_0</ID>786 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>240</ID>
<type>DE_OR8</type>
<position>51.5,-25.5</position>
<input>
<ID>IN_0</ID>297 </input>
<input>
<ID>IN_1</ID>296 </input>
<input>
<ID>IN_2</ID>270 </input>
<input>
<ID>IN_3</ID>253 </input>
<input>
<ID>IN_4</ID>250 </input>
<input>
<ID>IN_5</ID>250 </input>
<input>
<ID>IN_6</ID>251 </input>
<input>
<ID>IN_7</ID>252 </input>
<output>
<ID>OUT</ID>309 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>241</ID>
<type>DA_FROM</type>
<position>3,-19</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>242</ID>
<type>DA_FROM</type>
<position>3,-21</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>243</ID>
<type>DA_FROM</type>
<position>3,-24</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>574</ID>
<type>DA_FROM</type>
<position>149,-104</position>
<input>
<ID>IN_0</ID>796 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>244</ID>
<type>DA_FROM</type>
<position>3,-26</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp1</lparam></gate>
<gate>
<ID>245</ID>
<type>DA_FROM</type>
<position>3,-29</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>246</ID>
<type>DA_FROM</type>
<position>3,-31</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>569</ID>
<type>AA_AND2</type>
<position>169,-118</position>
<input>
<ID>IN_0</ID>803 </input>
<input>
<ID>IN_1</ID>804 </input>
<output>
<ID>OUT</ID>790 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>247</ID>
<type>AE_SMALL_INVERTER</type>
<position>11.5,-31</position>
<input>
<ID>IN_0</ID>303 </input>
<output>
<ID>OUT_0</ID>304 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>248</ID>
<type>DA_FROM</type>
<position>3,-34</position>
<input>
<ID>IN_0</ID>305 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>3,-36</position>
<input>
<ID>IN_0</ID>306 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>250</ID>
<type>DA_FROM</type>
<position>3,-41</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>251</ID>
<type>DE_TO</type>
<position>59.5,-25.5</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1in</lparam></gate>
<gate>
<ID>252</ID>
<type>DA_FROM</type>
<position>3,-16</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add1</lparam></gate>
<gate>
<ID>512</ID>
<type>DA_FROM</type>
<position>3,-122</position>
<input>
<ID>IN_0</ID>755 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>305</ID>
<type>AA_AND2</type>
<position>96,-40</position>
<input>
<ID>IN_0</ID>519 </input>
<input>
<ID>IN_1</ID>520 </input>
<output>
<ID>OUT</ID>503 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>DA_FROM</type>
<position>76,-39</position>
<input>
<ID>IN_0</ID>519 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>308</ID>
<type>AA_AND2</type>
<position>96,-10</position>
<input>
<ID>IN_0</ID>490 </input>
<input>
<ID>IN_1</ID>489 </input>
<output>
<ID>OUT</ID>509 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>516</ID>
<type>AA_AND2</type>
<position>23,-103</position>
<input>
<ID>IN_0</ID>747 </input>
<input>
<ID>IN_1</ID>746 </input>
<output>
<ID>OUT</ID>743 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>309</ID>
<type>AA_AND2</type>
<position>81.5,-11</position>
<input>
<ID>IN_0</ID>500 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>489 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>658</ID>
<type>DA_FROM</type>
<position>149,-136</position>
<input>
<ID>IN_0</ID>887 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>311</ID>
<type>DA_FROM</type>
<position>76,-7</position>
<input>
<ID>IN_0</ID>490 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_AND2</type>
<position>96,-25</position>
<input>
<ID>IN_0</ID>512 </input>
<input>
<ID>IN_1</ID>513 </input>
<output>
<ID>OUT</ID>506 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>520</ID>
<type>AA_AND2</type>
<position>23,-118</position>
<input>
<ID>IN_0</ID>753 </input>
<input>
<ID>IN_1</ID>754 </input>
<output>
<ID>OUT</ID>740 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>313</ID>
<type>AA_AND2</type>
<position>96,-30</position>
<input>
<ID>IN_0</ID>514 </input>
<input>
<ID>IN_1</ID>516 </input>
<output>
<ID>OUT</ID>505 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>315</ID>
<type>DA_FROM</type>
<position>76,-10</position>
<input>
<ID>IN_0</ID>500 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>316</ID>
<type>DA_FROM</type>
<position>76,-12</position>
<input>
<ID>IN_0</ID>501 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>524</ID>
<type>DE_OR8</type>
<position>51.5,-108.5</position>
<input>
<ID>IN_0</ID>745 </input>
<input>
<ID>IN_1</ID>744 </input>
<input>
<ID>IN_2</ID>743 </input>
<input>
<ID>IN_3</ID>742 </input>
<input>
<ID>IN_4</ID>739 </input>
<input>
<ID>IN_5</ID>739 </input>
<input>
<ID>IN_6</ID>740 </input>
<input>
<ID>IN_7</ID>741 </input>
<output>
<ID>OUT</ID>757 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>317</ID>
<type>DA_FROM</type>
<position>76,-14</position>
<input>
<ID>IN_0</ID>502 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>318</ID>
<type>DE_OR8</type>
<position>124.5,-25.5</position>
<input>
<ID>IN_0</ID>509 </input>
<input>
<ID>IN_1</ID>508 </input>
<input>
<ID>IN_2</ID>507 </input>
<input>
<ID>IN_3</ID>506 </input>
<input>
<ID>IN_4</ID>503 </input>
<input>
<ID>IN_5</ID>503 </input>
<input>
<ID>IN_6</ID>504 </input>
<input>
<ID>IN_7</ID>505 </input>
<output>
<ID>OUT</ID>521 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>666</ID>
<type>DA_FROM</type>
<position>149,-158</position>
<input>
<ID>IN_0</ID>903 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>319</ID>
<type>DA_FROM</type>
<position>76,-19</position>
<input>
<ID>IN_0</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>625</ID>
<type>DA_FROM</type>
<position>76,-163</position>
<input>
<ID>IN_0</ID>880 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>320</ID>
<type>DA_FROM</type>
<position>76,-21</position>
<input>
<ID>IN_0</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>656</ID>
<type>AA_AND2</type>
<position>169,-159</position>
<input>
<ID>IN_0</ID>903 </input>
<input>
<ID>IN_1</ID>904 </input>
<output>
<ID>OUT</ID>890 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>321</ID>
<type>DA_FROM</type>
<position>76,-24</position>
<input>
<ID>IN_0</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>322</ID>
<type>DA_FROM</type>
<position>76,-26</position>
<input>
<ID>IN_0</ID>513 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp2</lparam></gate>
<gate>
<ID>323</ID>
<type>DA_FROM</type>
<position>76,-29</position>
<input>
<ID>IN_0</ID>514 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>629</ID>
<type>AA_AND2</type>
<position>96,-149</position>
<input>
<ID>IN_0</ID>873 </input>
<input>
<ID>IN_1</ID>874 </input>
<output>
<ID>OUT</ID>867 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>324</ID>
<type>DA_FROM</type>
<position>76,-31</position>
<input>
<ID>IN_0</ID>515 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>660</ID>
<type>DA_FROM</type>
<position>149,-143</position>
<input>
<ID>IN_0</ID>897 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>325</ID>
<type>AE_SMALL_INVERTER</type>
<position>84.5,-31</position>
<input>
<ID>IN_0</ID>515 </input>
<output>
<ID>OUT_0</ID>516 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>326</ID>
<type>DA_FROM</type>
<position>76,-34</position>
<input>
<ID>IN_0</ID>517 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>327</ID>
<type>DA_FROM</type>
<position>76,-36</position>
<input>
<ID>IN_0</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>633</ID>
<type>DA_FROM</type>
<position>76,-138</position>
<input>
<ID>IN_0</ID>863 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>328</ID>
<type>DA_FROM</type>
<position>76,-41</position>
<input>
<ID>IN_0</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>664</ID>
<type>DA_FROM</type>
<position>149,-153</position>
<input>
<ID>IN_0</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>329</ID>
<type>DE_TO</type>
<position>132.5,-25.5</position>
<input>
<ID>IN_0</ID>521 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2in</lparam></gate>
<gate>
<ID>330</ID>
<type>DA_FROM</type>
<position>76,-16</position>
<input>
<ID>IN_0</ID>522 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add2</lparam></gate>
<gate>
<ID>331</ID>
<type>AA_AND2</type>
<position>169,-40</position>
<input>
<ID>IN_0</ID>544 </input>
<input>
<ID>IN_1</ID>545 </input>
<output>
<ID>OUT</ID>528 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>637</ID>
<type>DA_FROM</type>
<position>76,-148</position>
<input>
<ID>IN_0</ID>873 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>332</ID>
<type>AA_AND2</type>
<position>169,-15</position>
<input>
<ID>IN_0</ID>527 </input>
<input>
<ID>IN_1</ID>547 </input>
<output>
<ID>OUT</ID>533 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>668</ID>
<type>DE_TO</type>
<position>205.5,-149.5</position>
<input>
<ID>IN_0</ID>907 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15in</lparam></gate>
<gate>
<ID>333</ID>
<type>DA_FROM</type>
<position>149,-39</position>
<input>
<ID>IN_0</ID>544 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>334</ID>
<type>AA_AND2</type>
<position>169,-10</position>
<input>
<ID>IN_0</ID>524 </input>
<input>
<ID>IN_1</ID>523 </input>
<output>
<ID>OUT</ID>534 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>335</ID>
<type>AA_AND2</type>
<position>154.5,-11</position>
<input>
<ID>IN_0</ID>525 </input>
<input>
<ID>IN_1</ID>526 </input>
<output>
<ID>OUT</ID>523 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>513</ID>
<type>AA_AND2</type>
<position>23,-93</position>
<input>
<ID>IN_0</ID>735 </input>
<input>
<ID>IN_1</ID>734 </input>
<output>
<ID>OUT</ID>745 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>336</ID>
<type>AA_AND2</type>
<position>169,-20</position>
<input>
<ID>IN_0</ID>536 </input>
<input>
<ID>IN_1</ID>535 </input>
<output>
<ID>OUT</ID>532 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>672</ID>
<type>AA_LABEL</type>
<position>-49,70</position>
<gparam>LABEL_TEXT Checkpoint 2 - Brandon Aikman</gparam>
<gparam>TEXT_HEIGHT 2.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>337</ID>
<type>DA_FROM</type>
<position>149,-7</position>
<input>
<ID>IN_0</ID>524 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>338</ID>
<type>AA_AND2</type>
<position>169,-25</position>
<input>
<ID>IN_0</ID>537 </input>
<input>
<ID>IN_1</ID>538 </input>
<output>
<ID>OUT</ID>531 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>339</ID>
<type>AA_AND2</type>
<position>169,-30</position>
<input>
<ID>IN_0</ID>539 </input>
<input>
<ID>IN_1</ID>541 </input>
<output>
<ID>OUT</ID>530 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>517</ID>
<type>DA_FROM</type>
<position>3,-90</position>
<input>
<ID>IN_0</ID>735 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>340</ID>
<type>AA_AND2</type>
<position>169,-35</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>543 </input>
<output>
<ID>OUT</ID>529 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>DA_FROM</type>
<position>149,-10</position>
<input>
<ID>IN_0</ID>525 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>342</ID>
<type>DA_FROM</type>
<position>149,-12</position>
<input>
<ID>IN_0</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>343</ID>
<type>DA_FROM</type>
<position>149,-14</position>
<input>
<ID>IN_0</ID>527 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>345</ID>
<type>DA_FROM</type>
<position>149,-19</position>
<input>
<ID>IN_0</ID>536 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>346</ID>
<type>DA_FROM</type>
<position>149,-21</position>
<input>
<ID>IN_0</ID>535 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>347</ID>
<type>DA_FROM</type>
<position>149,-24</position>
<input>
<ID>IN_0</ID>537 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>525</ID>
<type>DA_FROM</type>
<position>3,-102</position>
<input>
<ID>IN_0</ID>747 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>348</ID>
<type>DA_FROM</type>
<position>149,-26</position>
<input>
<ID>IN_0</ID>538 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp3</lparam></gate>
<gate>
<ID>349</ID>
<type>DA_FROM</type>
<position>149,-29</position>
<input>
<ID>IN_0</ID>539 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>351</ID>
<type>AE_SMALL_INVERTER</type>
<position>157.5,-31</position>
<input>
<ID>IN_0</ID>540 </input>
<output>
<ID>OUT_0</ID>541 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>529</ID>
<type>DA_FROM</type>
<position>3,-112</position>
<input>
<ID>IN_0</ID>750 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>352</ID>
<type>DA_FROM</type>
<position>149,-34</position>
<input>
<ID>IN_0</ID>542 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>353</ID>
<type>DA_FROM</type>
<position>149,-36</position>
<input>
<ID>IN_0</ID>543 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>355</ID>
<type>DE_TO</type>
<position>205.5,-25.5</position>
<input>
<ID>IN_0</ID>546 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3in</lparam></gate>
<gate>
<ID>357</ID>
<type>AA_AND2</type>
<position>96,-61</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>654 </input>
<output>
<ID>OUT</ID>651 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>AA_AND2</type>
<position>-50,-56</position>
<input>
<ID>IN_0</ID>580 </input>
<input>
<ID>IN_1</ID>608 </input>
<output>
<ID>OUT</ID>594 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>AA_AND2</type>
<position>-50,-51</position>
<input>
<ID>IN_0</ID>549 </input>
<input>
<ID>IN_1</ID>548 </input>
<output>
<ID>OUT</ID>595 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>362</ID>
<type>AA_AND2</type>
<position>-64.5,-52</position>
<input>
<ID>IN_0</ID>550 </input>
<input>
<ID>IN_1</ID>567 </input>
<output>
<ID>OUT</ID>548 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>363</ID>
<type>AA_AND2</type>
<position>-50,-61</position>
<input>
<ID>IN_0</ID>597 </input>
<input>
<ID>IN_1</ID>596 </input>
<output>
<ID>OUT</ID>593 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>365</ID>
<type>AA_AND2</type>
<position>-50,-66</position>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>599 </input>
<output>
<ID>OUT</ID>592 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>367</ID>
<type>AA_AND2</type>
<position>-50,-76</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>604 </input>
<output>
<ID>OUT</ID>586 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>576</ID>
<type>DA_FROM</type>
<position>149,-109</position>
<input>
<ID>IN_0</ID>799 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp11</lparam></gate>
<gate>
<ID>369</ID>
<type>DA_FROM</type>
<position>-70,-53</position>
<input>
<ID>IN_0</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>371</ID>
<type>DE_OR8</type>
<position>-21.5,-66.5</position>
<input>
<ID>IN_0</ID>595 </input>
<input>
<ID>IN_1</ID>594 </input>
<input>
<ID>IN_2</ID>593 </input>
<input>
<ID>IN_3</ID>592 </input>
<input>
<ID>IN_4</ID>584 </input>
<input>
<ID>IN_5</ID>584 </input>
<input>
<ID>IN_6</ID>586 </input>
<input>
<ID>IN_7</ID>590 </input>
<output>
<ID>OUT</ID>607 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>580</ID>
<type>DA_FROM</type>
<position>149,-119</position>
<input>
<ID>IN_0</ID>804 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>373</ID>
<type>DA_FROM</type>
<position>-70,-62</position>
<input>
<ID>IN_0</ID>596 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>375</ID>
<type>DA_FROM</type>
<position>-70,-67</position>
<input>
<ID>IN_0</ID>599 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp4</lparam></gate>
<gate>
<ID>584</ID>
<type>AA_AND2</type>
<position>-50,-134</position>
<input>
<ID>IN_0</ID>810 </input>
<input>
<ID>IN_1</ID>809 </input>
<output>
<ID>OUT</ID>820 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>377</ID>
<type>DA_FROM</type>
<position>-70,-72</position>
<input>
<ID>IN_0</ID>601 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>379</ID>
<type>DA_FROM</type>
<position>-70,-75</position>
<input>
<ID>IN_0</ID>603 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>588</ID>
<type>AA_AND2</type>
<position>-50,-159</position>
<input>
<ID>IN_0</ID>828 </input>
<input>
<ID>IN_1</ID>829 </input>
<output>
<ID>OUT</ID>815 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>DA_FROM</type>
<position>-70,-82</position>
<input>
<ID>IN_0</ID>606 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>383</ID>
<type>AA_AND2</type>
<position>96,-56</position>
<input>
<ID>IN_0</ID>646 </input>
<input>
<ID>IN_1</ID>678 </input>
<output>
<ID>OUT</ID>652 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>384</ID>
<type>AA_AND2</type>
<position>96,-76</position>
<input>
<ID>IN_0</ID>673 </input>
<input>
<ID>IN_1</ID>674 </input>
<output>
<ID>OUT</ID>648 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>551</ID>
<type>DA_FROM</type>
<position>76,-109</position>
<input>
<ID>IN_0</ID>774 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp10</lparam></gate>
<gate>
<ID>386</ID>
<type>DA_FROM</type>
<position>149,-72</position>
<input>
<ID>IN_0</ID>701 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>387</ID>
<type>DE_OR8</type>
<position>197.5,-66.5</position>
<input>
<ID>IN_0</ID>690 </input>
<input>
<ID>IN_1</ID>689 </input>
<input>
<ID>IN_2</ID>688 </input>
<input>
<ID>IN_3</ID>687 </input>
<input>
<ID>IN_4</ID>684 </input>
<input>
<ID>IN_5</ID>684 </input>
<input>
<ID>IN_6</ID>685 </input>
<input>
<ID>IN_7</ID>686 </input>
<output>
<ID>OUT</ID>707 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>388</ID>
<type>DA_FROM</type>
<position>149,-82</position>
<input>
<ID>IN_0</ID>706 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>389</ID>
<type>DA_FROM</type>
<position>-70,-57</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add4</lparam></gate>
<gate>
<ID>539</ID>
<type>AA_AND2</type>
<position>96,-93</position>
<input>
<ID>IN_0</ID>760 </input>
<input>
<ID>IN_1</ID>759 </input>
<output>
<ID>OUT</ID>770 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>390</ID>
<type>AA_AND2</type>
<position>23,-81</position>
<input>
<ID>IN_0</ID>638 </input>
<input>
<ID>IN_1</ID>639 </input>
<output>
<ID>OUT</ID>622 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>391</ID>
<type>AA_AND2</type>
<position>23,-56</position>
<input>
<ID>IN_0</ID>621 </input>
<input>
<ID>IN_1</ID>641 </input>
<output>
<ID>OUT</ID>627 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>392</ID>
<type>DA_FROM</type>
<position>3,-80</position>
<input>
<ID>IN_0</ID>638 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>393</ID>
<type>AA_AND2</type>
<position>23,-51</position>
<input>
<ID>IN_0</ID>618 </input>
<input>
<ID>IN_1</ID>617 </input>
<output>
<ID>OUT</ID>628 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>559</ID>
<type>DA_FROM</type>
<position>76,-99</position>
<input>
<ID>IN_0</ID>783 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add10</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_AND2</type>
<position>8.5,-52</position>
<input>
<ID>IN_0</ID>619 </input>
<input>
<ID>IN_1</ID>620 </input>
<output>
<ID>OUT</ID>617 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>395</ID>
<type>AA_AND2</type>
<position>23,-61</position>
<input>
<ID>IN_0</ID>630 </input>
<input>
<ID>IN_1</ID>629 </input>
<output>
<ID>OUT</ID>626 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>396</ID>
<type>DA_FROM</type>
<position>3,-48</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>547</ID>
<type>DE_OR8</type>
<position>124.5,-108.5</position>
<input>
<ID>IN_0</ID>770 </input>
<input>
<ID>IN_1</ID>769 </input>
<input>
<ID>IN_2</ID>768 </input>
<input>
<ID>IN_3</ID>767 </input>
<input>
<ID>IN_4</ID>764 </input>
<input>
<ID>IN_5</ID>764 </input>
<input>
<ID>IN_6</ID>765 </input>
<input>
<ID>IN_7</ID>766 </input>
<output>
<ID>OUT</ID>782 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>398</ID>
<type>AA_AND2</type>
<position>23,-71</position>
<input>
<ID>IN_0</ID>633 </input>
<input>
<ID>IN_1</ID>635 </input>
<output>
<ID>OUT</ID>624 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>399</ID>
<type>AA_AND2</type>
<position>23,-76</position>
<input>
<ID>IN_0</ID>636 </input>
<input>
<ID>IN_1</ID>637 </input>
<output>
<ID>OUT</ID>623 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>577</ID>
<type>DA_FROM</type>
<position>149,-112</position>
<input>
<ID>IN_0</ID>800 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>400</ID>
<type>DA_FROM</type>
<position>3,-51</position>
<input>
<ID>IN_0</ID>619 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>401</ID>
<type>DA_FROM</type>
<position>3,-53</position>
<input>
<ID>IN_0</ID>620 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>567</ID>
<type>AA_AND2</type>
<position>169,-108</position>
<input>
<ID>IN_0</ID>798 </input>
<input>
<ID>IN_1</ID>799 </input>
<output>
<ID>OUT</ID>792 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>402</ID>
<type>DA_FROM</type>
<position>3,-55</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>403</ID>
<type>DE_OR8</type>
<position>51.5,-66.5</position>
<input>
<ID>IN_0</ID>628 </input>
<input>
<ID>IN_1</ID>627 </input>
<input>
<ID>IN_2</ID>626 </input>
<input>
<ID>IN_3</ID>625 </input>
<input>
<ID>IN_4</ID>622 </input>
<input>
<ID>IN_5</ID>622 </input>
<input>
<ID>IN_6</ID>623 </input>
<input>
<ID>IN_7</ID>624 </input>
<output>
<ID>OUT</ID>640 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>581</ID>
<type>DE_TO</type>
<position>205.5,-108.5</position>
<input>
<ID>IN_0</ID>807 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11in</lparam></gate>
<gate>
<ID>404</ID>
<type>DA_FROM</type>
<position>3,-60</position>
<input>
<ID>IN_0</ID>630 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>555</ID>
<type>DA_FROM</type>
<position>76,-117</position>
<input>
<ID>IN_0</ID>778 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>406</ID>
<type>DA_FROM</type>
<position>3,-65</position>
<input>
<ID>IN_0</ID>631 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>407</ID>
<type>DA_FROM</type>
<position>3,-67</position>
<input>
<ID>IN_0</ID>632 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp5</lparam></gate>
<gate>
<ID>585</ID>
<type>AA_AND2</type>
<position>-64.5,-135</position>
<input>
<ID>IN_0</ID>811 </input>
<input>
<ID>IN_1</ID>812 </input>
<output>
<ID>OUT</ID>809 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>408</ID>
<type>DA_FROM</type>
<position>3,-70</position>
<input>
<ID>IN_0</ID>633 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>575</ID>
<type>DA_FROM</type>
<position>149,-107</position>
<input>
<ID>IN_0</ID>798 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>410</ID>
<type>AE_SMALL_INVERTER</type>
<position>11.5,-72</position>
<input>
<ID>IN_0</ID>634 </input>
<output>
<ID>OUT_0</ID>635 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>411</ID>
<type>DA_FROM</type>
<position>3,-75</position>
<input>
<ID>IN_0</ID>636 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>589</ID>
<type>DA_FROM</type>
<position>-70,-136</position>
<input>
<ID>IN_0</ID>812 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>412</ID>
<type>DA_FROM</type>
<position>3,-77</position>
<input>
<ID>IN_0</ID>637 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>413</ID>
<type>DA_FROM</type>
<position>3,-82</position>
<input>
<ID>IN_0</ID>639 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>563</ID>
<type>AA_AND2</type>
<position>169,-93</position>
<input>
<ID>IN_0</ID>785 </input>
<input>
<ID>IN_1</ID>784 </input>
<output>
<ID>OUT</ID>795 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>414</ID>
<type>DE_TO</type>
<position>59.5,-66.5</position>
<input>
<ID>IN_0</ID>640 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5in</lparam></gate>
<gate>
<ID>593</ID>
<type>DA_FROM</type>
<position>-70,-155</position>
<input>
<ID>IN_0</ID>826 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>416</ID>
<type>AA_AND2</type>
<position>96,-81</position>
<input>
<ID>IN_0</ID>675 </input>
<input>
<ID>IN_1</ID>676 </input>
<output>
<ID>OUT</ID>647 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>417</ID>
<type>DA_FROM</type>
<position>76,-80</position>
<input>
<ID>IN_0</ID>675 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_AND2</type>
<position>96,-51</position>
<input>
<ID>IN_0</ID>643 </input>
<input>
<ID>IN_1</ID>642 </input>
<output>
<ID>OUT</ID>653 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>419</ID>
<type>AA_AND2</type>
<position>81.5,-52</position>
<input>
<ID>IN_0</ID>644 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>642 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>597</ID>
<type>AA_AND2</type>
<position>96,-159</position>
<input>
<ID>IN_0</ID>878 </input>
<input>
<ID>IN_1</ID>879 </input>
<output>
<ID>OUT</ID>865 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>420</ID>
<type>DA_FROM</type>
<position>76,-48</position>
<input>
<ID>IN_0</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>421</ID>
<type>AA_AND2</type>
<position>96,-66</position>
<input>
<ID>IN_0</ID>656 </input>
<input>
<ID>IN_1</ID>669 </input>
<output>
<ID>OUT</ID>650 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>571</ID>
<type>DA_FROM</type>
<position>149,-95</position>
<input>
<ID>IN_0</ID>787 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>422</ID>
<type>AA_AND2</type>
<position>96,-71</position>
<input>
<ID>IN_0</ID>670 </input>
<input>
<ID>IN_1</ID>672 </input>
<output>
<ID>OUT</ID>649 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>423</ID>
<type>DA_FROM</type>
<position>76,-51</position>
<input>
<ID>IN_0</ID>644 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>601</ID>
<type>DA_FROM</type>
<position>-70,-140</position>
<input>
<ID>IN_0</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add12</lparam></gate>
<gate>
<ID>424</ID>
<type>DA_FROM</type>
<position>76,-53</position>
<input>
<ID>IN_0</ID>645 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>425</ID>
<type>DA_FROM</type>
<position>76,-55</position>
<input>
<ID>IN_0</ID>646 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>426</ID>
<type>DE_OR8</type>
<position>124.5,-66.5</position>
<input>
<ID>IN_0</ID>653 </input>
<input>
<ID>IN_1</ID>652 </input>
<input>
<ID>IN_2</ID>651 </input>
<input>
<ID>IN_3</ID>650 </input>
<input>
<ID>IN_4</ID>647 </input>
<input>
<ID>IN_5</ID>647 </input>
<input>
<ID>IN_6</ID>648 </input>
<input>
<ID>IN_7</ID>649 </input>
<output>
<ID>OUT</ID>677 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>427</ID>
<type>DA_FROM</type>
<position>76,-60</position>
<input>
<ID>IN_0</ID>655 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>605</ID>
<type>AA_AND2</type>
<position>23,-134</position>
<input>
<ID>IN_0</ID>835 </input>
<input>
<ID>IN_1</ID>834 </input>
<output>
<ID>OUT</ID>845 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>428</ID>
<type>DA_FROM</type>
<position>76,-62</position>
<input>
<ID>IN_0</ID>654 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>429</ID>
<type>DA_FROM</type>
<position>76,-65</position>
<input>
<ID>IN_0</ID>656 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>430</ID>
<type>DA_FROM</type>
<position>76,-67</position>
<input>
<ID>IN_0</ID>669 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp6</lparam></gate>
<gate>
<ID>431</ID>
<type>DA_FROM</type>
<position>76,-70</position>
<input>
<ID>IN_0</ID>670 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>609</ID>
<type>AA_AND2</type>
<position>23,-154</position>
<input>
<ID>IN_0</ID>850 </input>
<input>
<ID>IN_1</ID>852 </input>
<output>
<ID>OUT</ID>841 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>432</ID>
<type>DA_FROM</type>
<position>76,-72</position>
<input>
<ID>IN_0</ID>671 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>640</ID>
<type>DA_FROM</type>
<position>76,-155</position>
<input>
<ID>IN_0</ID>876 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>433</ID>
<type>AE_SMALL_INVERTER</type>
<position>84.5,-72</position>
<input>
<ID>IN_0</ID>671 </input>
<output>
<ID>OUT_0</ID>672 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>434</ID>
<type>DA_FROM</type>
<position>76,-75</position>
<input>
<ID>IN_0</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>435</ID>
<type>DA_FROM</type>
<position>76,-77</position>
<input>
<ID>IN_0</ID>674 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>613</ID>
<type>DA_FROM</type>
<position>3,-138</position>
<input>
<ID>IN_0</ID>838 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>436</ID>
<type>DA_FROM</type>
<position>76,-82</position>
<input>
<ID>IN_0</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>644</ID>
<type>DA_FROM</type>
<position>76,-165</position>
<input>
<ID>IN_0</ID>881 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>437</ID>
<type>DE_TO</type>
<position>132.5,-66.5</position>
<input>
<ID>IN_0</ID>677 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6in</lparam></gate>
<gate>
<ID>438</ID>
<type>DA_FROM</type>
<position>76,-57</position>
<input>
<ID>IN_0</ID>678 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add6</lparam></gate>
<gate>
<ID>439</ID>
<type>AA_AND2</type>
<position>169,-81</position>
<input>
<ID>IN_0</ID>705 </input>
<input>
<ID>IN_1</ID>706 </input>
<output>
<ID>OUT</ID>684 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>617</ID>
<type>DA_FROM</type>
<position>3,-150</position>
<input>
<ID>IN_0</ID>849 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp13</lparam></gate>
<gate>
<ID>440</ID>
<type>AA_AND2</type>
<position>169,-56</position>
<input>
<ID>IN_0</ID>683 </input>
<input>
<ID>IN_1</ID>708 </input>
<output>
<ID>OUT</ID>689 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>648</ID>
<type>AA_AND2</type>
<position>169,-139</position>
<input>
<ID>IN_0</ID>888 </input>
<input>
<ID>IN_1</ID>908 </input>
<output>
<ID>OUT</ID>894 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>441</ID>
<type>DA_FROM</type>
<position>149,-80</position>
<input>
<ID>IN_0</ID>705 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>442</ID>
<type>AA_AND2</type>
<position>169,-51</position>
<input>
<ID>IN_0</ID>680 </input>
<input>
<ID>IN_1</ID>679 </input>
<output>
<ID>OUT</ID>690 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>443</ID>
<type>AA_AND2</type>
<position>154.5,-52</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>682 </input>
<output>
<ID>OUT</ID>679 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>621</ID>
<type>DA_FROM</type>
<position>3,-160</position>
<input>
<ID>IN_0</ID>854 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>444</ID>
<type>AA_AND2</type>
<position>169,-61</position>
<input>
<ID>IN_0</ID>692 </input>
<input>
<ID>IN_1</ID>691 </input>
<output>
<ID>OUT</ID>688 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>652</ID>
<type>AA_AND2</type>
<position>169,-144</position>
<input>
<ID>IN_0</ID>897 </input>
<input>
<ID>IN_1</ID>896 </input>
<output>
<ID>OUT</ID>893 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>445</ID>
<type>DA_FROM</type>
<position>149,-48</position>
<input>
<ID>IN_0</ID>680 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>446</ID>
<type>AA_AND2</type>
<position>169,-66</position>
<input>
<ID>IN_0</ID>698 </input>
<input>
<ID>IN_1</ID>699 </input>
<output>
<ID>OUT</ID>687 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>447</ID>
<type>AA_AND2</type>
<position>169,-71</position>
<input>
<ID>IN_0</ID>700 </input>
<input>
<ID>IN_1</ID>702 </input>
<output>
<ID>OUT</ID>686 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>448</ID>
<type>AA_AND2</type>
<position>169,-76</position>
<input>
<ID>IN_0</ID>703 </input>
<input>
<ID>IN_1</ID>704 </input>
<output>
<ID>OUT</ID>685 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>449</ID>
<type>DA_FROM</type>
<position>149,-51</position>
<input>
<ID>IN_0</ID>681 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>615</ID>
<type>DA_FROM</type>
<position>3,-143</position>
<input>
<ID>IN_0</ID>847 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>450</ID>
<type>DA_FROM</type>
<position>149,-53</position>
<input>
<ID>IN_0</ID>682 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>451</ID>
<type>DA_FROM</type>
<position>149,-55</position>
<input>
<ID>IN_0</ID>683 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>452</ID>
<type>DA_FROM</type>
<position>149,-60</position>
<input>
<ID>IN_0</ID>692 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>453</ID>
<type>DA_FROM</type>
<position>149,-62</position>
<input>
<ID>IN_0</ID>691 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>603</ID>
<type>AA_AND2</type>
<position>23,-139</position>
<input>
<ID>IN_0</ID>838 </input>
<input>
<ID>IN_1</ID>858 </input>
<output>
<ID>OUT</ID>844 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>454</ID>
<type>DA_FROM</type>
<position>149,-65</position>
<input>
<ID>IN_0</ID>698 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>455</ID>
<type>DA_FROM</type>
<position>149,-67</position>
<input>
<ID>IN_0</ID>699 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp7</lparam></gate>
<gate>
<ID>456</ID>
<type>DA_FROM</type>
<position>149,-70</position>
<input>
<ID>IN_0</ID>700 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>457</ID>
<type>AE_SMALL_INVERTER</type>
<position>157.5,-72</position>
<input>
<ID>IN_0</ID>701 </input>
<output>
<ID>OUT_0</ID>702 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>623</ID>
<type>DE_TO</type>
<position>59.5,-149.5</position>
<input>
<ID>IN_0</ID>857 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13in</lparam></gate>
<gate>
<ID>458</ID>
<type>DA_FROM</type>
<position>149,-75</position>
<input>
<ID>IN_0</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>459</ID>
<type>DA_FROM</type>
<position>149,-77</position>
<input>
<ID>IN_0</ID>704 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>460</ID>
<type>DE_TO</type>
<position>205.5,-66.5</position>
<input>
<ID>IN_0</ID>707 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7in</lparam></gate>
<gate>
<ID>461</ID>
<type>AA_AND2</type>
<position>96,-103</position>
<input>
<ID>IN_0</ID>772 </input>
<input>
<ID>IN_1</ID>771 </input>
<output>
<ID>OUT</ID>768 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>611</ID>
<type>DA_FROM</type>
<position>3,-134</position>
<input>
<ID>IN_0</ID>836 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>462</ID>
<type>AA_AND2</type>
<position>-50,-123</position>
<input>
<ID>IN_0</ID>730 </input>
<input>
<ID>IN_1</ID>731 </input>
<output>
<ID>OUT</ID>714 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>463</ID>
<type>AA_AND2</type>
<position>-50,-98</position>
<input>
<ID>IN_0</ID>713 </input>
<input>
<ID>IN_1</ID>733 </input>
<output>
<ID>OUT</ID>719 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>641</ID>
<type>AE_SMALL_INVERTER</type>
<position>84.5,-155</position>
<input>
<ID>IN_0</ID>876 </input>
<output>
<ID>OUT_0</ID>877 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>464</ID>
<type>DA_FROM</type>
<position>-70,-122</position>
<input>
<ID>IN_0</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>465</ID>
<type>AA_AND2</type>
<position>-50,-93</position>
<input>
<ID>IN_0</ID>710 </input>
<input>
<ID>IN_1</ID>709 </input>
<output>
<ID>OUT</ID>720 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>631</ID>
<type>DA_FROM</type>
<position>76,-134</position>
<input>
<ID>IN_0</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>466</ID>
<type>AA_AND2</type>
<position>-64.5,-94</position>
<input>
<ID>IN_0</ID>711 </input>
<input>
<ID>IN_1</ID>712 </input>
<output>
<ID>OUT</ID>709 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>467</ID>
<type>AA_AND2</type>
<position>-50,-103</position>
<input>
<ID>IN_0</ID>722 </input>
<input>
<ID>IN_1</ID>721 </input>
<output>
<ID>OUT</ID>718 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>645</ID>
<type>DE_TO</type>
<position>132.5,-149.5</position>
<input>
<ID>IN_0</ID>882 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14in</lparam></gate>
<gate>
<ID>468</ID>
<type>DA_FROM</type>
<position>-70,-90</position>
<input>
<ID>IN_0</ID>710 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>619</ID>
<type>AE_SMALL_INVERTER</type>
<position>11.5,-155</position>
<input>
<ID>IN_0</ID>851 </input>
<output>
<ID>OUT_0</ID>852 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>470</ID>
<type>DA_FROM</type>
<position>149,-140</position>
<input>
<ID>IN_0</ID>908 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add15</lparam></gate>
<gate>
<ID>649</ID>
<type>DA_FROM</type>
<position>149,-163</position>
<input>
<ID>IN_0</ID>905 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>472</ID>
<type>AA_AND2</type>
<position>-50,-118</position>
<input>
<ID>IN_0</ID>728 </input>
<input>
<ID>IN_1</ID>729 </input>
<output>
<ID>OUT</ID>715 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>473</ID>
<type>DA_FROM</type>
<position>-70,-93</position>
<input>
<ID>IN_0</ID>711 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>639</ID>
<type>DA_FROM</type>
<position>76,-153</position>
<input>
<ID>IN_0</ID>875 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>474</ID>
<type>AA_AND2</type>
<position>23,-149</position>
<input>
<ID>IN_0</ID>848 </input>
<input>
<ID>IN_1</ID>849 </input>
<output>
<ID>OUT</ID>842 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>475</ID>
<type>DA_FROM</type>
<position>-70,-95</position>
<input>
<ID>IN_0</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>653</ID>
<type>DA_FROM</type>
<position>149,-131</position>
<input>
<ID>IN_0</ID>885 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>476</ID>
<type>DA_FROM</type>
<position>-70,-97</position>
<input>
<ID>IN_0</ID>713 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>477</ID>
<type>DE_OR8</type>
<position>-21.5,-108.5</position>
<input>
<ID>IN_0</ID>720 </input>
<input>
<ID>IN_1</ID>719 </input>
<input>
<ID>IN_2</ID>718 </input>
<input>
<ID>IN_3</ID>717 </input>
<input>
<ID>IN_4</ID>714 </input>
<input>
<ID>IN_5</ID>714 </input>
<input>
<ID>IN_6</ID>715 </input>
<input>
<ID>IN_7</ID>716 </input>
<output>
<ID>OUT</ID>732 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>627</ID>
<type>AA_AND2</type>
<position>81.5,-135</position>
<input>
<ID>IN_0</ID>861 </input>
<input>
<ID>IN_1</ID>862 </input>
<output>
<ID>OUT</ID>859 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>478</ID>
<type>DA_FROM</type>
<position>3,-145</position>
<input>
<ID>IN_0</ID>846 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>479</ID>
<type>DA_FROM</type>
<position>-70,-102</position>
<input>
<ID>IN_0</ID>722 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>657</ID>
<type>DA_FROM</type>
<position>149,-134</position>
<input>
<ID>IN_0</ID>886 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>480</ID>
<type>DA_FROM</type>
<position>-70,-104</position>
<input>
<ID>IN_0</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>481</ID>
<type>DA_FROM</type>
<position>3,-140</position>
<input>
<ID>IN_0</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add13</lparam></gate>
<gate>
<ID>519</ID>
<type>AA_AND2</type>
<position>23,-113</position>
<input>
<ID>IN_0</ID>750 </input>
<input>
<ID>IN_1</ID>752 </input>
<output>
<ID>OUT</ID>741 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>482</ID>
<type>DA_FROM</type>
<position>-70,-107</position>
<input>
<ID>IN_0</ID>723 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>483</ID>
<type>DA_FROM</type>
<position>-70,-109</position>
<input>
<ID>IN_0</ID>724 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp8</lparam></gate>
<gate>
<ID>661</ID>
<type>DA_FROM</type>
<position>149,-145</position>
<input>
<ID>IN_0</ID>896 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>484</ID>
<type>DA_FROM</type>
<position>3,-155</position>
<input>
<ID>IN_0</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>485</ID>
<type>DA_FROM</type>
<position>-70,-112</position>
<input>
<ID>IN_0</ID>725 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>635</ID>
<type>DA_FROM</type>
<position>76,-143</position>
<input>
<ID>IN_0</ID>872 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>486</ID>
<type>DA_FROM</type>
<position>-70,-114</position>
<input>
<ID>IN_0</ID>726 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>487</ID>
<type>AE_SMALL_INVERTER</type>
<position>-61.5,-114</position>
<input>
<ID>IN_0</ID>726 </input>
<output>
<ID>OUT_0</ID>727 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>665</ID>
<type>AE_SMALL_INVERTER</type>
<position>157.5,-155</position>
<input>
<ID>IN_0</ID>901 </input>
<output>
<ID>OUT_0</ID>902 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>488</ID>
<type>DA_FROM</type>
<position>-70,-117</position>
<input>
<ID>IN_0</ID>728 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>489</ID>
<type>DA_FROM</type>
<position>-70,-119</position>
<input>
<ID>IN_0</ID>729 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>527</ID>
<type>DA_FROM</type>
<position>3,-107</position>
<input>
<ID>IN_0</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>490</ID>
<type>DA_FROM</type>
<position>-70,-124</position>
<input>
<ID>IN_0</ID>731 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>491</ID>
<type>DE_TO</type>
<position>-13.5,-108.5</position>
<input>
<ID>IN_0</ID>732 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8in</lparam></gate>
<gate>
<ID>492</ID>
<type>AA_AND2</type>
<position>96,-98</position>
<input>
<ID>IN_0</ID>763 </input>
<input>
<ID>IN_1</ID>783 </input>
<output>
<ID>OUT</ID>769 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>493</ID>
<type>AA_AND2</type>
<position>96,-118</position>
<input>
<ID>IN_0</ID>778 </input>
<input>
<ID>IN_1</ID>779 </input>
<output>
<ID>OUT</ID>765 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>515</ID>
<type>AA_AND2</type>
<position>8.5,-94</position>
<input>
<ID>IN_0</ID>736 </input>
<input>
<ID>IN_1</ID>737 </input>
<output>
<ID>OUT</ID>734 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>494</ID>
<type>DA_FROM</type>
<position>149,-99</position>
<input>
<ID>IN_0</ID>808 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add11</lparam></gate>
<gate>
<ID>495</ID>
<type>DA_FROM</type>
<position>149,-114</position>
<input>
<ID>IN_0</ID>801 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>496</ID>
<type>DE_OR8</type>
<position>197.5,-108.5</position>
<input>
<ID>IN_0</ID>795 </input>
<input>
<ID>IN_1</ID>794 </input>
<input>
<ID>IN_2</ID>793 </input>
<input>
<ID>IN_3</ID>792 </input>
<input>
<ID>IN_4</ID>789 </input>
<input>
<ID>IN_5</ID>789 </input>
<input>
<ID>IN_6</ID>790 </input>
<input>
<ID>IN_7</ID>791 </input>
<output>
<ID>OUT</ID>807 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>497</ID>
<type>DA_FROM</type>
<position>149,-124</position>
<input>
<ID>IN_0</ID>806 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>535</ID>
<type>DE_TO</type>
<position>59.5,-108.5</position>
<input>
<ID>IN_0</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9in</lparam></gate>
<gate>
<ID>498</ID>
<type>DA_FROM</type>
<position>-70,-131</position>
<input>
<ID>IN_0</ID>810 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>499</ID>
<type>AA_AND2</type>
<position>-50,-164</position>
<input>
<ID>IN_0</ID>830 </input>
<input>
<ID>IN_1</ID>831 </input>
<output>
<ID>OUT</ID>814 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>500</ID>
<type>DA_FROM</type>
<position>-70,-99</position>
<input>
<ID>IN_0</ID>733 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add8</lparam></gate>
<gate>
<ID>501</ID>
<type>DA_FROM</type>
<position>-70,-143</position>
<input>
<ID>IN_0</ID>822 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>523</ID>
<type>DA_FROM</type>
<position>3,-97</position>
<input>
<ID>IN_0</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>502</ID>
<type>AA_AND2</type>
<position>-50,-154</position>
<input>
<ID>IN_0</ID>825 </input>
<input>
<ID>IN_1</ID>827 </input>
<output>
<ID>OUT</ID>816 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>503</ID>
<type>DA_FROM</type>
<position>-70,-163</position>
<input>
<ID>IN_0</ID>830 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>504</ID>
<type>DA_FROM</type>
<position>-70,-138</position>
<input>
<ID>IN_0</ID>813 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>505</ID>
<type>DA_FROM</type>
<position>-70,-160</position>
<input>
<ID>IN_0</ID>829 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>543</ID>
<type>AA_AND2</type>
<position>96,-113</position>
<input>
<ID>IN_0</ID>775 </input>
<input>
<ID>IN_1</ID>777 </input>
<output>
<ID>OUT</ID>766 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>506</ID>
<type>DA_FROM</type>
<position>-70,-148</position>
<input>
<ID>IN_0</ID>823 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>508</ID>
<type>AE_SMALL_INVERTER</type>
<position>-61.5,-155</position>
<input>
<ID>IN_0</ID>826 </input>
<output>
<ID>OUT_0</ID>827 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>531</ID>
<type>AE_SMALL_INVERTER</type>
<position>11.5,-114</position>
<input>
<ID>IN_0</ID>751 </input>
<output>
<ID>OUT_0</ID>752 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>510</ID>
<type>AA_AND2</type>
<position>23,-98</position>
<input>
<ID>IN_0</ID>738 </input>
<input>
<ID>IN_1</ID>758 </input>
<output>
<ID>OUT</ID>744 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>511</ID>
<type>DE_TO</type>
<position>-13.5,-149.5</position>
<input>
<ID>IN_0</ID>832 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12in</lparam></gate>
<gate>
<ID>514</ID>
<type>DA_FROM</type>
<position>-70,-153</position>
<input>
<ID>IN_0</ID>825 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>518</ID>
<type>AA_AND2</type>
<position>23,-108</position>
<input>
<ID>IN_0</ID>748 </input>
<input>
<ID>IN_1</ID>749 </input>
<output>
<ID>OUT</ID>742 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>522</ID>
<type>DA_FROM</type>
<position>3,-95</position>
<input>
<ID>IN_0</ID>737 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>528</ID>
<type>DA_FROM</type>
<position>3,-109</position>
<input>
<ID>IN_0</ID>749 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp9</lparam></gate>
<gate>
<ID>532</ID>
<type>DA_FROM</type>
<position>3,-117</position>
<input>
<ID>IN_0</ID>753 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>536</ID>
<type>DA_FROM</type>
<position>3,-99</position>
<input>
<ID>IN_0</ID>758 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add9</lparam></gate>
<gate>
<ID>538</ID>
<type>DA_FROM</type>
<position>76,-122</position>
<input>
<ID>IN_0</ID>780 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>540</ID>
<type>AA_AND2</type>
<position>81.5,-94</position>
<input>
<ID>IN_0</ID>761 </input>
<input>
<ID>IN_1</ID>762 </input>
<output>
<ID>OUT</ID>759 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>544</ID>
<type>DA_FROM</type>
<position>76,-93</position>
<input>
<ID>IN_0</ID>761 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>548</ID>
<type>DA_FROM</type>
<position>76,-102</position>
<input>
<ID>IN_0</ID>772 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>552</ID>
<type>DA_FROM</type>
<position>76,-112</position>
<input>
<ID>IN_0</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>556</ID>
<type>DA_FROM</type>
<position>76,-119</position>
<input>
<ID>IN_0</ID>779 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>560</ID>
<type>AA_AND2</type>
<position>169,-123</position>
<input>
<ID>IN_0</ID>805 </input>
<input>
<ID>IN_1</ID>806 </input>
<output>
<ID>OUT</ID>789 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>564</ID>
<type>AA_AND2</type>
<position>154.5,-94</position>
<input>
<ID>IN_0</ID>786 </input>
<input>
<ID>IN_1</ID>787 </input>
<output>
<ID>OUT</ID>784 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>568</ID>
<type>AA_AND2</type>
<position>169,-113</position>
<input>
<ID>IN_0</ID>800 </input>
<input>
<ID>IN_1</ID>802 </input>
<output>
<ID>OUT</ID>791 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>572</ID>
<type>DA_FROM</type>
<position>149,-97</position>
<input>
<ID>IN_0</ID>788 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>578</ID>
<type>AE_SMALL_INVERTER</type>
<position>157.5,-114</position>
<input>
<ID>IN_0</ID>801 </input>
<output>
<ID>OUT_0</ID>802 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>579</ID>
<type>DA_FROM</type>
<position>149,-117</position>
<input>
<ID>IN_0</ID>803 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>582</ID>
<type>AA_AND2</type>
<position>96,-144</position>
<input>
<ID>IN_0</ID>872 </input>
<input>
<ID>IN_1</ID>871 </input>
<output>
<ID>OUT</ID>868 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>583</ID>
<type>AA_AND2</type>
<position>-50,-139</position>
<input>
<ID>IN_0</ID>813 </input>
<input>
<ID>IN_1</ID>833 </input>
<output>
<ID>OUT</ID>819 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>586</ID>
<type>AA_AND2</type>
<position>-50,-144</position>
<input>
<ID>IN_0</ID>822 </input>
<input>
<ID>IN_1</ID>821 </input>
<output>
<ID>OUT</ID>818 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>587</ID>
<type>AA_AND2</type>
<position>-50,-149</position>
<input>
<ID>IN_0</ID>823 </input>
<input>
<ID>IN_1</ID>824 </input>
<output>
<ID>OUT</ID>817 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>590</ID>
<type>DE_OR8</type>
<position>-21.5,-149.5</position>
<input>
<ID>IN_0</ID>820 </input>
<input>
<ID>IN_1</ID>819 </input>
<input>
<ID>IN_2</ID>818 </input>
<input>
<ID>IN_3</ID>817 </input>
<input>
<ID>IN_4</ID>814 </input>
<input>
<ID>IN_5</ID>814 </input>
<input>
<ID>IN_6</ID>815 </input>
<input>
<ID>IN_7</ID>816 </input>
<output>
<ID>OUT</ID>832 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>591</ID>
<type>DA_FROM</type>
<position>-70,-145</position>
<input>
<ID>IN_0</ID>821 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>592</ID>
<type>DA_FROM</type>
<position>-70,-150</position>
<input>
<ID>IN_0</ID>824 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp12</lparam></gate>
<gate>
<ID>594</ID>
<type>DA_FROM</type>
<position>-70,-158</position>
<input>
<ID>IN_0</ID>828 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>595</ID>
<type>DA_FROM</type>
<position>-70,-165</position>
<input>
<ID>IN_0</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>596</ID>
<type>AA_AND2</type>
<position>96,-139</position>
<input>
<ID>IN_0</ID>863 </input>
<input>
<ID>IN_1</ID>883 </input>
<output>
<ID>OUT</ID>869 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>598</ID>
<type>DA_FROM</type>
<position>149,-155</position>
<input>
<ID>IN_0</ID>901 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>599</ID>
<type>DE_OR8</type>
<position>197.5,-149.5</position>
<input>
<ID>IN_0</ID>895 </input>
<input>
<ID>IN_1</ID>894 </input>
<input>
<ID>IN_2</ID>893 </input>
<input>
<ID>IN_3</ID>892 </input>
<input>
<ID>IN_4</ID>889 </input>
<input>
<ID>IN_5</ID>889 </input>
<input>
<ID>IN_6</ID>890 </input>
<input>
<ID>IN_7</ID>891 </input>
<output>
<ID>OUT</ID>907 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>600</ID>
<type>DA_FROM</type>
<position>149,-165</position>
<input>
<ID>IN_0</ID>906 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>602</ID>
<type>AA_AND2</type>
<position>23,-164</position>
<input>
<ID>IN_0</ID>855 </input>
<input>
<ID>IN_1</ID>856 </input>
<output>
<ID>OUT</ID>839 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>604</ID>
<type>DA_FROM</type>
<position>3,-163</position>
<input>
<ID>IN_0</ID>855 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>606</ID>
<type>AA_AND2</type>
<position>8.5,-135</position>
<input>
<ID>IN_0</ID>836 </input>
<input>
<ID>IN_1</ID>837 </input>
<output>
<ID>OUT</ID>834 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>607</ID>
<type>AA_AND2</type>
<position>23,-144</position>
<input>
<ID>IN_0</ID>847 </input>
<input>
<ID>IN_1</ID>846 </input>
<output>
<ID>OUT</ID>843 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>608</ID>
<type>DA_FROM</type>
<position>3,-131</position>
<input>
<ID>IN_0</ID>835 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>610</ID>
<type>AA_AND2</type>
<position>23,-159</position>
<input>
<ID>IN_0</ID>853 </input>
<input>
<ID>IN_1</ID>854 </input>
<output>
<ID>OUT</ID>840 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>612</ID>
<type>DA_FROM</type>
<position>3,-136</position>
<input>
<ID>IN_0</ID>837 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>614</ID>
<type>DE_OR8</type>
<position>51.5,-149.5</position>
<input>
<ID>IN_0</ID>845 </input>
<input>
<ID>IN_1</ID>844 </input>
<input>
<ID>IN_2</ID>843 </input>
<input>
<ID>IN_3</ID>842 </input>
<input>
<ID>IN_4</ID>839 </input>
<input>
<ID>IN_5</ID>839 </input>
<input>
<ID>IN_6</ID>840 </input>
<input>
<ID>IN_7</ID>841 </input>
<output>
<ID>OUT</ID>857 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>616</ID>
<type>DA_FROM</type>
<position>3,-148</position>
<input>
<ID>IN_0</ID>848 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>618</ID>
<type>DA_FROM</type>
<position>3,-153</position>
<input>
<ID>IN_0</ID>850 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>620</ID>
<type>DA_FROM</type>
<position>3,-158</position>
<input>
<ID>IN_0</ID>853 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>622</ID>
<type>DA_FROM</type>
<position>3,-165</position>
<input>
<ID>IN_0</ID>856 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>624</ID>
<type>AA_AND2</type>
<position>96,-164</position>
<input>
<ID>IN_0</ID>880 </input>
<input>
<ID>IN_1</ID>881 </input>
<output>
<ID>OUT</ID>864 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>626</ID>
<type>AA_AND2</type>
<position>96,-134</position>
<input>
<ID>IN_0</ID>860 </input>
<input>
<ID>IN_1</ID>859 </input>
<output>
<ID>OUT</ID>870 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>628</ID>
<type>DA_FROM</type>
<position>76,-131</position>
<input>
<ID>IN_0</ID>860 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>630</ID>
<type>AA_AND2</type>
<position>96,-154</position>
<input>
<ID>IN_0</ID>875 </input>
<input>
<ID>IN_1</ID>877 </input>
<output>
<ID>OUT</ID>866 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>632</ID>
<type>DA_FROM</type>
<position>76,-136</position>
<input>
<ID>IN_0</ID>862 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>634</ID>
<type>DE_OR8</type>
<position>124.5,-149.5</position>
<input>
<ID>IN_0</ID>870 </input>
<input>
<ID>IN_1</ID>869 </input>
<input>
<ID>IN_2</ID>868 </input>
<input>
<ID>IN_3</ID>867 </input>
<input>
<ID>IN_4</ID>864 </input>
<input>
<ID>IN_5</ID>864 </input>
<input>
<ID>IN_6</ID>865 </input>
<input>
<ID>IN_7</ID>866 </input>
<output>
<ID>OUT</ID>882 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>636</ID>
<type>DA_FROM</type>
<position>76,-145</position>
<input>
<ID>IN_0</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>638</ID>
<type>DA_FROM</type>
<position>76,-150</position>
<input>
<ID>IN_0</ID>874 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp14</lparam></gate>
<gate>
<ID>642</ID>
<type>DA_FROM</type>
<position>76,-158</position>
<input>
<ID>IN_0</ID>878 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>643</ID>
<type>DA_FROM</type>
<position>76,-160</position>
<input>
<ID>IN_0</ID>879 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>646</ID>
<type>DA_FROM</type>
<position>76,-140</position>
<input>
<ID>IN_0</ID>883 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add14</lparam></gate>
<gate>
<ID>647</ID>
<type>AA_AND2</type>
<position>169,-164</position>
<input>
<ID>IN_0</ID>905 </input>
<input>
<ID>IN_1</ID>906 </input>
<output>
<ID>OUT</ID>889 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>650</ID>
<type>AA_AND2</type>
<position>169,-134</position>
<input>
<ID>IN_0</ID>885 </input>
<input>
<ID>IN_1</ID>884 </input>
<output>
<ID>OUT</ID>895 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>651</ID>
<type>AA_AND2</type>
<position>154.5,-135</position>
<input>
<ID>IN_0</ID>886 </input>
<input>
<ID>IN_1</ID>887 </input>
<output>
<ID>OUT</ID>884 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>654</ID>
<type>AA_AND2</type>
<position>169,-149</position>
<input>
<ID>IN_0</ID>898 </input>
<input>
<ID>IN_1</ID>899 </input>
<output>
<ID>OUT</ID>892 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>655</ID>
<type>AA_AND2</type>
<position>169,-154</position>
<input>
<ID>IN_0</ID>900 </input>
<input>
<ID>IN_1</ID>902 </input>
<output>
<ID>OUT</ID>891 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>659</ID>
<type>DA_FROM</type>
<position>149,-138</position>
<input>
<ID>IN_0</ID>888 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>662</ID>
<type>DA_FROM</type>
<position>149,-148</position>
<input>
<ID>IN_0</ID>898 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>663</ID>
<type>DA_FROM</type>
<position>149,-150</position>
<input>
<ID>IN_0</ID>899 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inp15</lparam></gate>
<gate>
<ID>667</ID>
<type>DA_FROM</type>
<position>149,-160</position>
<input>
<ID>IN_0</ID>904 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>671</ID>
<type>AA_LABEL</type>
<position>-57.5,76.5</position>
<gparam>LABEL_TEXT Mano Machine</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>888 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-138,166,-138</points>
<connection>
<GID>659</GID>
<name>IN_0</name></connection>
<connection>
<GID>648</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>743 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-107,37,-103</points>
<intersection>-107 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-107,48.5,-107</points>
<connection>
<GID>524</GID>
<name>IN_2</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-103,37,-103</points>
<connection>
<GID>516</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>41 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-25,-24.5,-25</points>
<connection>
<GID>45</GID>
<name>IN_3</name></connection>
<connection>
<GID>23</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>129 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,15,16,16.5</points>
<intersection>15 2</intersection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,16.5,16,16.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,15,17.5,15</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>65 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,46,64,50.5</points>
<intersection>46 2</intersection>
<intersection>50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,50.5,64,50.5</points>
<connection>
<GID>110</GID>
<name>OUT_2</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64,46,65,46</points>
<connection>
<GID>104</GID>
<name>IN_6</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>848 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-148,20,-148</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<connection>
<GID>474</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-61.5,-11,-53,-11</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<connection>
<GID>5</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>728 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-117,-53,-117</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<connection>
<GID>472</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-9,-62,-7</points>
<intersection>-9 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-9,-53,-9</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-68,-7,-62,-7</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>35 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-10,-67.5,-10</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<connection>
<GID>9</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>36 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-12,-67.5,-12</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<connection>
<GID>9</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>884 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157.5,-135,166,-135</points>
<connection>
<GID>651</GID>
<name>OUT</name></connection>
<connection>
<GID>650</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>723 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-107,-53,-107</points>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<connection>
<GID>469</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>37 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-14,-53,-14</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<connection>
<GID>21</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>732 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-108.5,-15.5,-108.5</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<intersection>-17.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-17.5,-108.5,-17.5,-108.5</points>
<connection>
<GID>477</GID>
<name>OUT</name></connection>
<intersection>-108.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>38 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-40,-34,-28</points>
<intersection>-40 2</intersection>
<intersection>-29 1</intersection>
<intersection>-28 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-29,-24.5,-29</points>
<connection>
<GID>45</GID>
<name>IN_4</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-40,-34,-40</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-34,-28,-24.5,-28</points>
<connection>
<GID>45</GID>
<name>IN_5</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>898 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-148,166,-148</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<connection>
<GID>654</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>39 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-35,-35,-27</points>
<intersection>-35 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,-27,-24.5,-27</points>
<connection>
<GID>45</GID>
<name>IN_6</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-35,-35,-35</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>40 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-30,-36,-26</points>
<intersection>-30 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-26,-24.5,-26</points>
<connection>
<GID>45</GID>
<name>IN_7</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-30,-36,-30</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>736 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-93,5.5,-93</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>5.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5.5,-93,5.5,-93</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>42 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-24,-36,-20</points>
<intersection>-24 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-24,-24.5,-24</points>
<connection>
<GID>45</GID>
<name>IN_2</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-20,-36,-20</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>43 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-23,-35,-15</points>
<intersection>-23 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-15,-35,-15</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-35,-23,-24.5,-23</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>44 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-22,-34,-10</points>
<intersection>-22 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-22,-24.5,-22</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-10,-34,-10</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>892 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-149,194.5,-149</points>
<connection>
<GID>654</GID>
<name>OUT</name></connection>
<connection>
<GID>599</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>731 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-124,-53,-124</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<connection>
<GID>462</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>45 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-21,-53,-21</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>22</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>740 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-118,38,-110</points>
<intersection>-118 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-110,48.5,-110</points>
<connection>
<GID>524</GID>
<name>IN_6</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-118,38,-118</points>
<connection>
<GID>520</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>46 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-19,-53,-19</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>906 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-165,166,-165</points>
<connection>
<GID>600</GID>
<name>IN_0</name></connection>
<connection>
<GID>647</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>47 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-24,-53,-24</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<connection>
<GID>23</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>48 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-26,-53,-26</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<connection>
<GID>23</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>768 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-107,110,-103</points>
<intersection>-107 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-107,121.5,-107</points>
<connection>
<GID>547</GID>
<name>IN_2</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-103,110,-103</points>
<connection>
<GID>461</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>751 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-114,9.5,-114</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>9.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>9.5,-114,9.5,-114</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<intersection>-114 1</intersection></vsegment></shape></wire>
<wire>
<ID>49 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-29,-53,-29</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>51 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-31,-63.5,-31</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<connection>
<GID>51</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>52 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-31,-53,-31</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>772 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-102,93,-102</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<connection>
<GID>461</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>739 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-123,39,-111</points>
<intersection>-123 2</intersection>
<intersection>-112 1</intersection>
<intersection>-111 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-112,48.5,-112</points>
<connection>
<GID>524</GID>
<name>IN_4</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-123,39,-123</points>
<connection>
<GID>509</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>39,-111,48.5,-111</points>
<connection>
<GID>524</GID>
<name>IN_5</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>53 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-34,-53,-34</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>748 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-107,20,-107</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<connection>
<GID>518</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>54 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-36,-53,-36</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>55 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-39,-53,-39</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>56 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-41,-53,-41</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>776 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>78,-114,82.5,-114</points>
<connection>
<GID>553</GID>
<name>IN_0</name></connection>
<intersection>82.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>82.5,-114,82.5,-114</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>-114 3</intersection></vsegment></shape></wire>
<wire>
<ID>759 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-94,93,-94</points>
<connection>
<GID>540</GID>
<name>OUT</name></connection>
<connection>
<GID>539</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>57 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,34.5,65,40</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>61.5,34.5,65,34.5</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>752 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-114,20,-114</points>
<connection>
<GID>531</GID>
<name>OUT_0</name></connection>
<connection>
<GID>519</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>58 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,36.5,64,41</points>
<intersection>36.5 2</intersection>
<intersection>41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,41,65,41</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,36.5,64,36.5</points>
<connection>
<GID>123</GID>
<name>OUT_1</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>59 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,38.5,63,42</points>
<intersection>38.5 2</intersection>
<intersection>42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,42,65,42</points>
<connection>
<GID>104</GID>
<name>IN_2</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,38.5,63,38.5</points>
<connection>
<GID>123</GID>
<name>OUT_2</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>60 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,40.5,62,43</points>
<intersection>40.5 2</intersection>
<intersection>43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,43,65,43</points>
<connection>
<GID>104</GID>
<name>IN_3</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,40.5,62,40.5</points>
<connection>
<GID>123</GID>
<name>OUT_3</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>127 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,31,17.5,31</points>
<connection>
<GID>148</GID>
<name>IN_2</name></connection>
<intersection>16 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>16,30.5,16,31</points>
<intersection>30.5 5</intersection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>15,30.5,16,30.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>16 4</intersection></hsegment></shape></wire>
<wire>
<ID>63 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,44,62,46.5</points>
<intersection>44 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,44,65,44</points>
<connection>
<GID>104</GID>
<name>IN_4</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,46.5,62,46.5</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>128 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,28.5,16,30</points>
<intersection>28.5 1</intersection>
<intersection>30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,28.5,16,28.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,30,17.5,30</points>
<connection>
<GID>148</GID>
<name>IN_3</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>881 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-165,93,-165</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<connection>
<GID>624</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>64 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,45,63,48.5</points>
<intersection>45 1</intersection>
<intersection>48.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,45,65,45</points>
<connection>
<GID>104</GID>
<name>IN_5</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,48.5,63,48.5</points>
<connection>
<GID>110</GID>
<name>OUT_1</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>807 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>201.5,-108.5,203.5,-108.5</points>
<connection>
<GID>581</GID>
<name>IN_0</name></connection>
<intersection>201.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>201.5,-108.5,201.5,-108.5</points>
<connection>
<GID>496</GID>
<name>OUT</name></connection>
<intersection>-108.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>130 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,12.5,16,12.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>16 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>16,12.5,16,13</points>
<intersection>12.5 1</intersection>
<intersection>13 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>16,13,17.5,13</points>
<connection>
<GID>149</GID>
<name>IN_2</name></connection>
<intersection>16 2</intersection></hsegment></shape></wire>
<wire>
<ID>66 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,47,65,52.5</points>
<connection>
<GID>104</GID>
<name>IN_7</name></connection>
<intersection>52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,52.5,65,52.5</points>
<connection>
<GID>110</GID>
<name>OUT_3</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>131 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,10.5,16,12</points>
<intersection>10.5 2</intersection>
<intersection>12 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>15,10.5,16,10.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>16,12,17.5,12</points>
<connection>
<GID>149</GID>
<name>IN_3</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>67 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,30,68,38</points>
<connection>
<GID>104</GID>
<name>clock</name></connection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,30,68,30</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>132 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,14.5,16,14.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>16 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>16,14,16,14.5</points>
<intersection>14 7</intersection>
<intersection>14.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>16,14,17.5,14</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>16 6</intersection></hsegment></shape></wire>
<wire>
<ID>885 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-133,157,-131</points>
<intersection>-133 1</intersection>
<intersection>-131 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-133,166,-133</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-131,157,-131</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment></shape></wire>
<wire>
<ID>68 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,47,77,47</points>
<connection>
<GID>104</GID>
<name>OUT_7</name></connection>
<connection>
<GID>135</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>133 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,76,16.5,79</points>
<intersection>76 1</intersection>
<intersection>79 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,76,17.5,76</points>
<connection>
<GID>151</GID>
<name>IN_B_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,79,16.5,79</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,46,84.5,46</points>
<connection>
<GID>104</GID>
<name>OUT_6</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>795 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-105,185,-93</points>
<intersection>-105 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-105,194.5,-105</points>
<connection>
<GID>496</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-93,185,-93</points>
<connection>
<GID>563</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>134 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,75,16,77</points>
<intersection>75 2</intersection>
<intersection>77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,77,16,77</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,75,17.5,75</points>
<connection>
<GID>151</GID>
<name>IN_B_1</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>70 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,45,77,45</points>
<connection>
<GID>104</GID>
<name>OUT_5</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>71 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,44,84.5,44</points>
<connection>
<GID>104</GID>
<name>OUT_4</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>889 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-164,185,-152</points>
<intersection>-164 2</intersection>
<intersection>-153 1</intersection>
<intersection>-152 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-153,194.5,-153</points>
<connection>
<GID>599</GID>
<name>IN_4</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-164,185,-164</points>
<connection>
<GID>647</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>185,-152,194.5,-152</points>
<connection>
<GID>599</GID>
<name>IN_5</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>72 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,43,77,43</points>
<connection>
<GID>104</GID>
<name>OUT_3</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>73 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,42,84.5,42</points>
<connection>
<GID>104</GID>
<name>OUT_2</name></connection>
<connection>
<GID>142</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,41,77,41</points>
<connection>
<GID>104</GID>
<name>OUT_1</name></connection>
<connection>
<GID>143</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,40,84.5,40</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<connection>
<GID>144</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>893 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-148,183,-144</points>
<intersection>-148 1</intersection>
<intersection>-144 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183,-148,194.5,-148</points>
<connection>
<GID>599</GID>
<name>IN_2</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-144,183,-144</points>
<connection>
<GID>652</GID>
<name>OUT</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>76 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-25.5,-15.5,-25.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<connection>
<GID>45</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>77 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,25,20.5,27</points>
<connection>
<GID>149</GID>
<name>carry_in</name></connection>
<connection>
<GID>148</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>78 </ID>
<shape>
<vsegment>
<ID>12</ID>
<points>20.5,61,20.5,63</points>
<connection>
<GID>150</GID>
<name>carry_in</name></connection>
<connection>
<GID>151</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>79 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,43,20.5,45</points>
<connection>
<GID>150</GID>
<name>carry_out</name></connection>
<connection>
<GID>148</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>769 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-106,111,-98</points>
<intersection>-106 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-98,111,-98</points>
<connection>
<GID>492</GID>
<name>OUT</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111,-106,121.5,-106</points>
<connection>
<GID>547</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>80 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,3,31.5,3</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>81 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,3,20.5,9</points>
<connection>
<GID>149</GID>
<name>carry_out</name></connection>
<intersection>3 1</intersection>
<intersection>5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,3,25,3</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>20.5,5,31.5,5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,79,26.5,80</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>20.5,79,20.5,80</points>
<connection>
<GID>151</GID>
<name>carry_in</name></connection>
<intersection>80 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>20.5,80,26.5,80</points>
<intersection>20.5 1</intersection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,69,16,70.5</points>
<intersection>69 4</intersection>
<intersection>70.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>15,70.5,16,70.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>16,69,17.5,69</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>773 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-107,93,-107</points>
<connection>
<GID>550</GID>
<name>IN_0</name></connection>
<connection>
<GID>542</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>84 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,68.5,16,68.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,68,16,68.5</points>
<intersection>68 4</intersection>
<intersection>68.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>16,68,17.5,68</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<intersection>16 3</intersection></hsegment></shape></wire>
<wire>
<ID>85 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,67,17.5,67</points>
<connection>
<GID>151</GID>
<name>IN_2</name></connection>
<intersection>16 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>16,66.5,16,67</points>
<intersection>66.5 5</intersection>
<intersection>67 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>15,66.5,16,66.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>16 4</intersection></hsegment></shape></wire>
<wire>
<ID>86 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,64.5,16,66</points>
<intersection>64.5 1</intersection>
<intersection>66 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,64.5,16,64.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,66,17.5,66</points>
<connection>
<GID>151</GID>
<name>IN_3</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>87 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,51,16,52.5</points>
<intersection>51 2</intersection>
<intersection>52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,52.5,16,52.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,51,17.5,51</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>777 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-114,93,-114</points>
<connection>
<GID>554</GID>
<name>OUT_0</name></connection>
<connection>
<GID>543</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>88 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,48.5,16,49</points>
<intersection>48.5 1</intersection>
<intersection>49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,48.5,16,48.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,49,17.5,49</points>
<connection>
<GID>150</GID>
<name>IN_2</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>89 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,46.5,16,48</points>
<intersection>46.5 1</intersection>
<intersection>48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,46.5,16,46.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,48,17.5,48</points>
<connection>
<GID>150</GID>
<name>IN_3</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>90 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,50,16,50.5</points>
<intersection>50 1</intersection>
<intersection>50.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,50,17.5,50</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,50.5,16,50.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>91 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,33,16,34.5</points>
<intersection>33 2</intersection>
<intersection>34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,34.5,16,34.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,33,17.5,33</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>781 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-124,93,-124</points>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<connection>
<GID>537</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>92 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,32.5,16,32.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>16 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>16,32,16,32.5</points>
<intersection>32 5</intersection>
<intersection>32.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>16,32,17.5,32</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>16 4</intersection></hsegment></shape></wire>
<wire>
<ID>135 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,74,15.5,75</points>
<intersection>74 1</intersection>
<intersection>75 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,74,17.5,74</points>
<connection>
<GID>151</GID>
<name>IN_B_2</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,75,15.5,75</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,73,17.5,73</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<connection>
<GID>151</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>137 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,55,17.5,55</points>
<connection>
<GID>150</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>197</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>815 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-159,-35,-151</points>
<intersection>-159 2</intersection>
<intersection>-151 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,-151,-24.5,-151</points>
<connection>
<GID>590</GID>
<name>IN_6</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-159,-35,-159</points>
<connection>
<GID>588</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>138 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,56,15.5,57</points>
<intersection>56 2</intersection>
<intersection>57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,57,15.5,57</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,56,17.5,56</points>
<connection>
<GID>150</GID>
<name>IN_B_2</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>300 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-24,20,-24</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<connection>
<GID>234</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>139 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,57,16,59</points>
<intersection>57 2</intersection>
<intersection>59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,59,16,59</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,57,17.5,57</points>
<connection>
<GID>150</GID>
<name>IN_B_1</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>140 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,58,16.5,61</points>
<intersection>58 1</intersection>
<intersection>61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,58,17.5,58</points>
<connection>
<GID>150</GID>
<name>IN_B_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,61,16.5,61</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,37,17.5,37</points>
<connection>
<GID>148</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>201</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>803 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-117,166,-117</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<connection>
<GID>569</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>142 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,38,15.5,39</points>
<intersection>38 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,39,15.5,39</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,38,17.5,38</points>
<connection>
<GID>148</GID>
<name>IN_B_2</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,39,16,41</points>
<intersection>39 2</intersection>
<intersection>41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,41,16,41</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,39,17.5,39</points>
<connection>
<GID>148</GID>
<name>IN_B_1</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>883 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-140,93,-140</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-140,93,-140</points>
<connection>
<GID>596</GID>
<name>IN_1</name></connection>
<intersection>-140 1</intersection></vsegment></shape></wire>
<wire>
<ID>222 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,40,16.5,43</points>
<intersection>40 1</intersection>
<intersection>43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,40,17.5,40</points>
<connection>
<GID>148</GID>
<name>IN_B_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,43,16.5,43</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>545 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-41,166,-41</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>223 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,19,17.5,19</points>
<connection>
<GID>149</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>205</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>224 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,20,15.5,21</points>
<intersection>20 2</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,21,15.5,21</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,20,17.5,20</points>
<connection>
<GID>149</GID>
<name>IN_B_2</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>225 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,21,16,23</points>
<intersection>21 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,23,16,23</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,21,17.5,21</points>
<connection>
<GID>149</GID>
<name>IN_B_1</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>775 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-112,93,-112</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<connection>
<GID>543</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>226 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,22,16.5,25</points>
<intersection>22 2</intersection>
<intersection>25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,25,16.5,25</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,22,17.5,22</points>
<connection>
<GID>149</GID>
<name>IN_B_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>227 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-16,-53,-16</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<connection>
<GID>21</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>228 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>27,72,28,72</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>27 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>27,71.5,27,72</points>
<intersection>71.5 7</intersection>
<intersection>72 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>25.5,71.5,27,71.5</points>
<connection>
<GID>151</GID>
<name>OUT_1</name></connection>
<intersection>27 6</intersection></hsegment></shape></wire>
<wire>
<ID>891 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-154,183,-150</points>
<intersection>-154 2</intersection>
<intersection>-150 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183,-150,194.5,-150</points>
<connection>
<GID>599</GID>
<name>IN_7</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-154,183,-154</points>
<connection>
<GID>655</GID>
<name>OUT</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>230 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,70,28,70</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,70,27,70.5</points>
<intersection>70 1</intersection>
<intersection>70.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>25.5,70.5,27,70.5</points>
<connection>
<GID>151</GID>
<name>OUT_2</name></connection>
<intersection>27 3</intersection></hsegment></shape></wire>
<wire>
<ID>231 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,72.5,27,74</points>
<intersection>72.5 2</intersection>
<intersection>74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,74,28,74</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,72.5,27,72.5</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>232 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,68,27,69.5</points>
<intersection>68 1</intersection>
<intersection>69.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,68,28,68</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,69.5,27,69.5</points>
<connection>
<GID>151</GID>
<name>OUT_3</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>233 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,54.5,27,56</points>
<intersection>54.5 2</intersection>
<intersection>56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,56,28,56</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,54.5,27,54.5</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>783 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-99,93,-99</points>
<connection>
<GID>559</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-99,93,-99</points>
<connection>
<GID>492</GID>
<name>IN_1</name></connection>
<intersection>-99 1</intersection></vsegment></shape></wire>
<wire>
<ID>234 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,53.5,27,54</points>
<intersection>53.5 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,53.5,27,53.5</points>
<connection>
<GID>150</GID>
<name>OUT_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,54,28,54</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>235 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,52.5,27,52.5</points>
<connection>
<GID>150</GID>
<name>OUT_2</name></connection>
<intersection>27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,52,27,52.5</points>
<intersection>52 4</intersection>
<intersection>52.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>27,52,28,52</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>27 3</intersection></hsegment></shape></wire>
<wire>
<ID>236 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,50,27,51.5</points>
<intersection>50 1</intersection>
<intersection>51.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,50,28,50</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,51.5,27,51.5</points>
<connection>
<GID>150</GID>
<name>OUT_3</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>237 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,36.5,27,38</points>
<intersection>36.5 2</intersection>
<intersection>38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,38,28,38</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,36.5,27,36.5</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>771 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-104,93,-104</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-104,93,-104</points>
<connection>
<GID>461</GID>
<name>IN_1</name></connection>
<intersection>-104 1</intersection></vsegment></shape></wire>
<wire>
<ID>238 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,35.5,27,35.5</points>
<connection>
<GID>148</GID>
<name>OUT_1</name></connection>
<intersection>27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,35.5,27,36</points>
<intersection>35.5 1</intersection>
<intersection>36 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>27,36,28,36</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>27 3</intersection></hsegment></shape></wire>
<wire>
<ID>239 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,34,27,34.5</points>
<intersection>34 1</intersection>
<intersection>34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,34,28,34</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,34.5,27,34.5</points>
<connection>
<GID>148</GID>
<name>OUT_2</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>240 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,32,27,33.5</points>
<intersection>32 1</intersection>
<intersection>33.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,32,28,32</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,33.5,27,33.5</points>
<connection>
<GID>148</GID>
<name>OUT_3</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>241 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,18,28,18</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>27 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>27,17.5,27,18</points>
<intersection>17.5 5</intersection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>25.5,17.5,27,17.5</points>
<connection>
<GID>149</GID>
<name>OUT_1</name></connection>
<intersection>27 4</intersection></hsegment></shape></wire>
<wire>
<ID>791 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-113,183,-109</points>
<intersection>-113 2</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183,-109,194.5,-109</points>
<connection>
<GID>496</GID>
<name>IN_7</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-113,183,-113</points>
<connection>
<GID>568</GID>
<name>OUT</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>242 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,16,27,16.5</points>
<intersection>16 1</intersection>
<intersection>16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,16,28,16</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,16.5,27,16.5</points>
<connection>
<GID>149</GID>
<name>OUT_2</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>243 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,18.5,27,20</points>
<intersection>18.5 1</intersection>
<intersection>20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,18.5,27,18.5</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,20,28,20</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>244 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,14,27,15.5</points>
<intersection>14 1</intersection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,14,28,14</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,15.5,27,15.5</points>
<connection>
<GID>149</GID>
<name>OUT_3</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>270 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-24,37,-20</points>
<intersection>-24 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-24,48.5,-24</points>
<connection>
<GID>240</GID>
<name>IN_2</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-20,37,-20</points>
<connection>
<GID>232</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>245 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-11,20,-11</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<connection>
<GID>230</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>779 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-119,93,-119</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-119,93,-119</points>
<connection>
<GID>493</GID>
<name>IN_1</name></connection>
<intersection>-119 1</intersection></vsegment></shape></wire>
<wire>
<ID>246 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-9,11,-7</points>
<intersection>-9 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-9,20,-9</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-7,11,-7</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>247 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-10,5.5,-10</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>5.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5.5,-10,5.5,-10</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>-10 1</intersection></vsegment></shape></wire>
<wire>
<ID>248 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-12,5.5,-12</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>5.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5.5,-12,5.5,-12</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>249 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-14,20,-14</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<connection>
<GID>228</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>799 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-109,166,-109</points>
<connection>
<GID>576</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-109,166,-109</points>
<connection>
<GID>567</GID>
<name>IN_1</name></connection>
<intersection>-109 1</intersection></vsegment></shape></wire>
<wire>
<ID>250 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-40,39,-28</points>
<intersection>-40 2</intersection>
<intersection>-29 1</intersection>
<intersection>-28 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-29,48.5,-29</points>
<connection>
<GID>240</GID>
<name>IN_4</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-40,39,-40</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>39,-28,48.5,-28</points>
<connection>
<GID>240</GID>
<name>IN_5</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>251 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-35,38,-27</points>
<intersection>-35 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-27,48.5,-27</points>
<connection>
<GID>240</GID>
<name>IN_6</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-35,38,-35</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>252 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-30,37,-26</points>
<intersection>-30 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-26,48.5,-26</points>
<connection>
<GID>240</GID>
<name>IN_7</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-30,37,-30</points>
<connection>
<GID>235</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>253 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-25,48.5,-25</points>
<connection>
<GID>240</GID>
<name>IN_3</name></connection>
<connection>
<GID>234</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>296 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-23,38,-15</points>
<intersection>-23 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-15,38,-15</points>
<connection>
<GID>228</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-23,48.5,-23</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>632 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-67,20,-67</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>20 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>20,-67,20,-67</points>
<connection>
<GID>397</GID>
<name>IN_1</name></connection>
<intersection>-67 1</intersection></vsegment></shape></wire>
<wire>
<ID>297 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-22,39,-10</points>
<intersection>-22 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-22,48.5,-22</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-10,39,-10</points>
<connection>
<GID>230</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>298 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-21,20,-21</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-21,20,-21</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>299 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-19,20,-19</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>636 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-75,20,-75</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<connection>
<GID>399</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>301 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-26,20,-26</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-26,20,-26</points>
<connection>
<GID>234</GID>
<name>IN_1</name></connection>
<intersection>-26 1</intersection></vsegment></shape></wire>
<wire>
<ID>302 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-29,20,-29</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<connection>
<GID>235</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>650 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99,-66,121.5,-66</points>
<connection>
<GID>426</GID>
<name>IN_3</name></connection>
<connection>
<GID>421</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>303 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-31,9.5,-31</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>9.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>9.5,-31,9.5,-31</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>-31 1</intersection></vsegment></shape></wire>
<wire>
<ID>304 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-31,20,-31</points>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection>
<connection>
<GID>235</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>512 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-24,93,-24</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<connection>
<GID>312</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>305 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-34,20,-34</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<connection>
<GID>236</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>306 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-36,20,-36</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-36,20,-36</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>-36 1</intersection></vsegment></shape></wire>
<wire>
<ID>670 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-70,93,-70</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<connection>
<GID>422</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>307 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-39,20,-39</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<connection>
<GID>227</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>308 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-41,20,-41</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<connection>
<GID>227</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>516 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-31,93,-31</points>
<connection>
<GID>325</GID>
<name>OUT_0</name></connection>
<connection>
<GID>313</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>309 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-25.5,57.5,-25.5</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>55.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>55.5,-25.5,55.5,-25.5</points>
<connection>
<GID>240</GID>
<name>OUT</name></connection>
<intersection>-25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>310 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-16,20,-16</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-16,20,-16</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>-16 1</intersection></vsegment></shape></wire>
<wire>
<ID>489 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-11,93,-11</points>
<connection>
<GID>309</GID>
<name>OUT</name></connection>
<connection>
<GID>308</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>527 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-14,166,-14</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<connection>
<GID>332</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>490 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-9,84,-7</points>
<intersection>-9 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-9,93,-9</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-7,84,-7</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>830 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-163,-53,-163</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<connection>
<GID>499</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>677 </ID>
<shape>
<hsegment>
<ID>11</ID>
<points>128.5,-66.5,130.5,-66.5</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<intersection>128.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>128.5,-66.5,128.5,-66.5</points>
<connection>
<GID>426</GID>
<name>OUT</name></connection>
<intersection>-66.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>500 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-10,78.5,-10</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-10,78.5,-10</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>-10 1</intersection></vsegment></shape></wire>
<wire>
<ID>708 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-57,166,-57</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>166 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>166,-57,166,-57</points>
<connection>
<GID>440</GID>
<name>IN_1</name></connection>
<intersection>-57 1</intersection></vsegment></shape></wire>
<wire>
<ID>501 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-12,78.5,-12</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-12,78.5,-12</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>523 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157.5,-11,166,-11</points>
<connection>
<GID>335</GID>
<name>OUT</name></connection>
<connection>
<GID>334</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>502 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-14,93,-14</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<connection>
<GID>306</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>825 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-153,-53,-153</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<connection>
<GID>502</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>503 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-40,112,-28</points>
<intersection>-40 2</intersection>
<intersection>-29 1</intersection>
<intersection>-28 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-29,121.5,-29</points>
<connection>
<GID>318</GID>
<name>IN_4</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-40,112,-40</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>112,-28,121.5,-28</points>
<connection>
<GID>318</GID>
<name>IN_5</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>681 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-51,151.5,-51</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>151.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>151.5,-51,151.5,-51</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>-51 1</intersection></vsegment></shape></wire>
<wire>
<ID>504 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-35,111,-27</points>
<intersection>-35 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-27,121.5,-27</points>
<connection>
<GID>318</GID>
<name>IN_6</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-35,111,-35</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>712 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-95,-67.5,-95</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>-67.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-67.5,-95,-67.5,-95</points>
<connection>
<GID>466</GID>
<name>IN_1</name></connection>
<intersection>-95 1</intersection></vsegment></shape></wire>
<wire>
<ID>505 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-30,110,-26</points>
<intersection>-30 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-26,121.5,-26</points>
<connection>
<GID>318</GID>
<name>IN_7</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-30,110,-30</points>
<connection>
<GID>313</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>543 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-36,166,-36</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-36,166,-36</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>-36 1</intersection></vsegment></shape></wire>
<wire>
<ID>506 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99,-25,121.5,-25</points>
<connection>
<GID>312</GID>
<name>OUT</name></connection>
<connection>
<GID>318</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>507 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-24,110,-20</points>
<intersection>-24 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-24,121.5,-24</points>
<connection>
<GID>318</GID>
<name>IN_2</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-20,110,-20</points>
<connection>
<GID>310</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>685 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-76,184,-68</points>
<intersection>-76 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-68,194.5,-68</points>
<connection>
<GID>387</GID>
<name>IN_6</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-76,184,-76</points>
<connection>
<GID>448</GID>
<name>OUT</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>508 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-23,111,-15</points>
<intersection>-23 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-15,111,-15</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111,-23,121.5,-23</points>
<connection>
<GID>318</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>716 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-113,-36,-109</points>
<intersection>-113 2</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-109,-24.5,-109</points>
<connection>
<GID>477</GID>
<name>IN_7</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-113,-36,-113</points>
<connection>
<GID>471</GID>
<name>OUT</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>509 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-22,112,-10</points>
<intersection>-22 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-22,121.5,-22</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-10,112,-10</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>531 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-25,194.5,-25</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<connection>
<GID>344</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>510 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-21,93,-21</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-21,93,-21</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>511 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-19,93,-19</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<connection>
<GID>310</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>513 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-26,93,-26</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-26,93,-26</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<intersection>-26 1</intersection></vsegment></shape></wire>
<wire>
<ID>514 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-29,93,-29</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<connection>
<GID>313</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>515 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>78,-31,82.5,-31</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>82.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>82.5,-31,82.5,-31</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>-31 3</intersection></vsegment></shape></wire>
<wire>
<ID>517 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-34,93,-34</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<connection>
<GID>314</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>518 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-36,93,-36</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-36,93,-36</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>-36 1</intersection></vsegment></shape></wire>
<wire>
<ID>519 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-39,93,-39</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<connection>
<GID>305</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>520 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-41,93,-41</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<connection>
<GID>305</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>521 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>128.5,-25.5,130.5,-25.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>128.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128.5,-25.5,128.5,-25.5</points>
<connection>
<GID>318</GID>
<name>OUT</name></connection>
<intersection>-25.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>522 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-16,93,-16</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-16,93,-16</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<intersection>-16 1</intersection></vsegment></shape></wire>
<wire>
<ID>524 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-9,157,-7</points>
<intersection>-9 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-9,166,-9</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-7,157,-7</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment></shape></wire>
<wire>
<ID>525 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-10,151.5,-10</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>151.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>151.5,-10,151.5,-10</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>-10 1</intersection></vsegment></shape></wire>
<wire>
<ID>526 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-12,151.5,-12</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>151.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>151.5,-12,151.5,-12</points>
<connection>
<GID>335</GID>
<name>IN_1</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>528 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-40,185,-28</points>
<intersection>-40 2</intersection>
<intersection>-29 1</intersection>
<intersection>-28 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-29,194.5,-29</points>
<connection>
<GID>344</GID>
<name>IN_4</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-40,185,-40</points>
<connection>
<GID>331</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>185,-28,194.5,-28</points>
<connection>
<GID>344</GID>
<name>IN_5</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>529 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-35,184,-27</points>
<intersection>-35 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-27,194.5,-27</points>
<connection>
<GID>344</GID>
<name>IN_6</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-35,184,-35</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>530 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-30,183,-26</points>
<intersection>-30 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183,-26,194.5,-26</points>
<connection>
<GID>344</GID>
<name>IN_7</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-30,183,-30</points>
<connection>
<GID>339</GID>
<name>OUT</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>532 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-24,183,-20</points>
<intersection>-24 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183,-24,194.5,-24</points>
<connection>
<GID>344</GID>
<name>IN_2</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-20,183,-20</points>
<connection>
<GID>336</GID>
<name>OUT</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>533 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-23,184,-15</points>
<intersection>-23 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172,-15,184,-15</points>
<connection>
<GID>332</GID>
<name>OUT</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184,-23,194.5,-23</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>534 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-22,185,-10</points>
<intersection>-22 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-22,194.5,-22</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-10,185,-10</points>
<connection>
<GID>334</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>535 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-21,166,-21</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-21,166,-21</points>
<connection>
<GID>336</GID>
<name>IN_1</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>903 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-158,166,-158</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<connection>
<GID>656</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>536 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-19,166,-19</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<connection>
<GID>336</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>537 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-24,166,-24</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<connection>
<GID>338</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>897 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-143,166,-143</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<connection>
<GID>652</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>538 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-26,166,-26</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-26,166,-26</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>-26 1</intersection></vsegment></shape></wire>
<wire>
<ID>539 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-29,166,-29</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<connection>
<GID>339</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>540 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>151,-31,155.5,-31</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>155.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>155.5,-31,155.5,-31</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>-31 3</intersection></vsegment></shape></wire>
<wire>
<ID>541 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>159.5,-31,166,-31</points>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection>
<connection>
<GID>339</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>901 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>151,-155,155.5,-155</points>
<connection>
<GID>598</GID>
<name>IN_0</name></connection>
<intersection>155.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>155.5,-155,155.5,-155</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>-155 3</intersection></vsegment></shape></wire>
<wire>
<ID>542 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-34,166,-34</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<connection>
<GID>340</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>544 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-39,166,-39</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>905 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-163,166,-163</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<connection>
<GID>647</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>546 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>201.5,-25.5,203.5,-25.5</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>201.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>201.5,-25.5,201.5,-25.5</points>
<connection>
<GID>344</GID>
<name>OUT</name></connection>
<intersection>-25.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>547 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-16,166,-16</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-16,166,-16</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<intersection>-16 1</intersection></vsegment></shape></wire>
<wire>
<ID>899 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-150,166,-150</points>
<connection>
<GID>663</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-150,166,-150</points>
<connection>
<GID>654</GID>
<name>IN_1</name></connection>
<intersection>-150 1</intersection></vsegment></shape></wire>
<wire>
<ID>548 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-61.5,-52,-53,-52</points>
<connection>
<GID>362</GID>
<name>OUT</name></connection>
<connection>
<GID>361</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>549 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-50,-62,-48</points>
<intersection>-50 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-50,-53,-50</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-68,-48,-62,-48</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>550 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-68,-51,-67.5,-51</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<intersection>-67.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-67.5,-51,-67.5,-51</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>-51 3</intersection></vsegment></shape></wire>
<wire>
<ID>567 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-53,-67.5,-53</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>-67.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-67.5,-53,-67.5,-53</points>
<connection>
<GID>362</GID>
<name>IN_1</name></connection>
<intersection>-53 1</intersection></vsegment></shape></wire>
<wire>
<ID>580 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-55,-53,-55</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<connection>
<GID>370</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>584 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-81,-34,-69</points>
<intersection>-81 2</intersection>
<intersection>-70 1</intersection>
<intersection>-69 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-70,-24.5,-70</points>
<connection>
<GID>371</GID>
<name>IN_4</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-81,-34,-81</points>
<connection>
<GID>358</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-34,-69,-24.5,-69</points>
<connection>
<GID>371</GID>
<name>IN_5</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>586 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-76,-35,-68</points>
<intersection>-76 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,-68,-24.5,-68</points>
<connection>
<GID>371</GID>
<name>IN_6</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-76,-35,-76</points>
<connection>
<GID>367</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>590 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-71,-36,-67</points>
<intersection>-71 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-67,-24.5,-67</points>
<connection>
<GID>371</GID>
<name>IN_7</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-71,-36,-71</points>
<connection>
<GID>366</GID>
<name>OUT</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>592 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-66,-24.5,-66</points>
<connection>
<GID>371</GID>
<name>IN_3</name></connection>
<connection>
<GID>365</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>593 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-65,-36,-61</points>
<intersection>-65 1</intersection>
<intersection>-61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-65,-24.5,-65</points>
<connection>
<GID>371</GID>
<name>IN_2</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-61,-36,-61</points>
<connection>
<GID>363</GID>
<name>OUT</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>594 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-64,-35,-56</points>
<intersection>-64 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-56,-35,-56</points>
<connection>
<GID>359</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-35,-64,-24.5,-64</points>
<connection>
<GID>371</GID>
<name>IN_1</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>595 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-63,-34,-51</points>
<intersection>-63 1</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-63,-24.5,-63</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-51,-34,-51</points>
<connection>
<GID>361</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>596 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-62,-53,-62</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>-53 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-53,-62,-53,-62</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<intersection>-62 1</intersection></vsegment></shape></wire>
<wire>
<ID>597 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-60,-53,-60</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<connection>
<GID>372</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>598 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-65,-53,-65</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<connection>
<GID>374</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>599 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-67,-53,-67</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>-53 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-53,-67,-53,-67</points>
<connection>
<GID>365</GID>
<name>IN_1</name></connection>
<intersection>-67 1</intersection></vsegment></shape></wire>
<wire>
<ID>600 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-70,-53,-70</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<connection>
<GID>366</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>601 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-72,-63.5,-72</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>-63.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-63.5,-72,-63.5,-72</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>-72 1</intersection></vsegment></shape></wire>
<wire>
<ID>602 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-72,-53,-72</points>
<connection>
<GID>378</GID>
<name>OUT_0</name></connection>
<connection>
<GID>366</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>603 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-75,-53,-75</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>604 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-77,-53,-77</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>-53 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-53,-77,-53,-77</points>
<connection>
<GID>367</GID>
<name>IN_1</name></connection>
<intersection>-77 1</intersection></vsegment></shape></wire>
<wire>
<ID>605 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-80,-53,-80</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<connection>
<GID>358</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>606 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-82,-53,-82</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<connection>
<GID>358</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>607 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-66.5,-15.5,-66.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>-17.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-17.5,-66.5,-17.5,-66.5</points>
<connection>
<GID>371</GID>
<name>OUT</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>608 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-57,-53,-57</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>-53 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-53,-57,-53,-57</points>
<connection>
<GID>359</GID>
<name>IN_1</name></connection>
<intersection>-57 1</intersection></vsegment></shape></wire>
<wire>
<ID>617 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-52,20,-52</points>
<connection>
<GID>394</GID>
<name>OUT</name></connection>
<connection>
<GID>393</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>618 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-50,11,-48</points>
<intersection>-50 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-50,20,-50</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-48,11,-48</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>619 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-51,5.5,-51</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>5.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>5.5,-51,5.5,-51</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>-51 1</intersection></vsegment></shape></wire>
<wire>
<ID>620 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-53,5.5,-53</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<intersection>5.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>5.5,-53,5.5,-53</points>
<connection>
<GID>394</GID>
<name>IN_1</name></connection>
<intersection>-53 1</intersection></vsegment></shape></wire>
<wire>
<ID>621 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-55,20,-55</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<connection>
<GID>391</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>622 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-81,39,-69</points>
<intersection>-81 2</intersection>
<intersection>-70 1</intersection>
<intersection>-69 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-70,48.5,-70</points>
<connection>
<GID>403</GID>
<name>IN_4</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-81,39,-81</points>
<connection>
<GID>390</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>39,-69,48.5,-69</points>
<connection>
<GID>403</GID>
<name>IN_5</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>623 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-76,38,-68</points>
<intersection>-76 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-68,48.5,-68</points>
<connection>
<GID>403</GID>
<name>IN_6</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-76,38,-76</points>
<connection>
<GID>399</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>624 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-71,37,-67</points>
<intersection>-71 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-67,48.5,-67</points>
<connection>
<GID>403</GID>
<name>IN_7</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-71,37,-71</points>
<connection>
<GID>398</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>625 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-66,48.5,-66</points>
<connection>
<GID>403</GID>
<name>IN_3</name></connection>
<connection>
<GID>397</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>626 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-65,37,-61</points>
<intersection>-65 1</intersection>
<intersection>-61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-65,48.5,-65</points>
<connection>
<GID>403</GID>
<name>IN_2</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-61,37,-61</points>
<connection>
<GID>395</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>627 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-64,38,-56</points>
<intersection>-64 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-56,38,-56</points>
<connection>
<GID>391</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-64,48.5,-64</points>
<connection>
<GID>403</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>628 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-63,39,-51</points>
<intersection>-63 1</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-63,48.5,-63</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-51,39,-51</points>
<connection>
<GID>393</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>629 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-62,20,-62</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>20 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>20,-62,20,-62</points>
<connection>
<GID>395</GID>
<name>IN_1</name></connection>
<intersection>-62 1</intersection></vsegment></shape></wire>
<wire>
<ID>630 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-60,20,-60</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<connection>
<GID>395</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>631 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-65,20,-65</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<connection>
<GID>397</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>633 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-70,20,-70</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<connection>
<GID>398</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>634 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-72,9.5,-72</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>9.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>9.5,-72,9.5,-72</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>-72 1</intersection></vsegment></shape></wire>
<wire>
<ID>635 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-72,20,-72</points>
<connection>
<GID>410</GID>
<name>OUT_0</name></connection>
<connection>
<GID>398</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>637 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-77,20,-77</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>20 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>20,-77,20,-77</points>
<connection>
<GID>399</GID>
<name>IN_1</name></connection>
<intersection>-77 1</intersection></vsegment></shape></wire>
<wire>
<ID>638 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-80,20,-80</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<connection>
<GID>390</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>639 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-82,20,-82</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<connection>
<GID>390</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>640 </ID>
<shape>
<hsegment>
<ID>9</ID>
<points>55.5,-66.5,57.5,-66.5</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>55.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>55.5,-66.5,55.5,-66.5</points>
<connection>
<GID>403</GID>
<name>OUT</name></connection>
<intersection>-66.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>794 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-106,184,-98</points>
<intersection>-106 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172,-98,184,-98</points>
<connection>
<GID>561</GID>
<name>OUT</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184,-106,194.5,-106</points>
<connection>
<GID>496</GID>
<name>IN_1</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>641 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-57,20,-57</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>20 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>20,-57,20,-57</points>
<connection>
<GID>391</GID>
<name>IN_1</name></connection>
<intersection>-57 1</intersection></vsegment></shape></wire>
<wire>
<ID>642 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-52,93,-52</points>
<connection>
<GID>419</GID>
<name>OUT</name></connection>
<connection>
<GID>418</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>804 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-119,166,-119</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-119,166,-119</points>
<connection>
<GID>569</GID>
<name>IN_1</name></connection>
<intersection>-119 1</intersection></vsegment></shape></wire>
<wire>
<ID>643 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-50,84,-48</points>
<intersection>-50 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-50,93,-50</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-48,84,-48</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>644 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-51,78.5,-51</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<intersection>78.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>78.5,-51,78.5,-51</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>-51 1</intersection></vsegment></shape></wire>
<wire>
<ID>798 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-107,166,-107</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<connection>
<GID>567</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>645 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-53,78.5,-53</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<connection>
<GID>419</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>646 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-55,93,-55</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<connection>
<GID>383</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>792 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-108,194.5,-108</points>
<connection>
<GID>567</GID>
<name>OUT</name></connection>
<connection>
<GID>496</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>647 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-81,112,-69</points>
<intersection>-81 2</intersection>
<intersection>-70 1</intersection>
<intersection>-69 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-70,121.5,-70</points>
<connection>
<GID>426</GID>
<name>IN_4</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-81,112,-81</points>
<connection>
<GID>416</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>112,-69,121.5,-69</points>
<connection>
<GID>426</GID>
<name>IN_5</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>648 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-76,111,-68</points>
<intersection>-76 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-68,121.5,-68</points>
<connection>
<GID>426</GID>
<name>IN_6</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-76,111,-76</points>
<connection>
<GID>384</GID>
<name>OUT</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>802 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>159.5,-114,166,-114</points>
<connection>
<GID>578</GID>
<name>OUT_0</name></connection>
<connection>
<GID>568</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>649 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-71,110,-67</points>
<intersection>-71 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-67,121.5,-67</points>
<connection>
<GID>426</GID>
<name>IN_7</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-71,110,-71</points>
<connection>
<GID>422</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>812 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-136,-67.5,-136</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<intersection>-67.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-67.5,-136,-67.5,-136</points>
<connection>
<GID>585</GID>
<name>IN_1</name></connection>
<intersection>-136 1</intersection></vsegment></shape></wire>
<wire>
<ID>651 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-65,110,-61</points>
<intersection>-65 1</intersection>
<intersection>-61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-65,121.5,-65</points>
<connection>
<GID>426</GID>
<name>IN_2</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-61,110,-61</points>
<connection>
<GID>357</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>652 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-64,111,-56</points>
<intersection>-64 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-56,111,-56</points>
<connection>
<GID>383</GID>
<name>OUT</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111,-64,121.5,-64</points>
<connection>
<GID>426</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>806 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-124,166,-124</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<connection>
<GID>560</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>653 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-63,112,-51</points>
<intersection>-63 1</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-63,121.5,-63</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-51,112,-51</points>
<connection>
<GID>418</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>654 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-62,93,-62</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>93 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>93,-62,93,-62</points>
<connection>
<GID>357</GID>
<name>IN_1</name></connection>
<intersection>-62 1</intersection></vsegment></shape></wire>
<wire>
<ID>800 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-112,166,-112</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<connection>
<GID>568</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>655 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-60,93,-60</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<connection>
<GID>357</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>656 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-65,93,-65</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<connection>
<GID>421</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>822 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-143,-53,-143</points>
<connection>
<GID>501</GID>
<name>IN_0</name></connection>
<connection>
<GID>586</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>669 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-67,93,-67</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>93 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>93,-67,93,-67</points>
<connection>
<GID>421</GID>
<name>IN_1</name></connection>
<intersection>-67 1</intersection></vsegment></shape></wire>
<wire>
<ID>816 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-154,-36,-150</points>
<intersection>-154 2</intersection>
<intersection>-150 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-150,-24.5,-150</points>
<connection>
<GID>590</GID>
<name>IN_7</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-154,-36,-154</points>
<connection>
<GID>502</GID>
<name>OUT</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>671 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>78,-72,82.5,-72</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<intersection>82.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>82.5,-72,82.5,-72</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>-72 3</intersection></vsegment></shape></wire>
<wire>
<ID>672 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-72,93,-72</points>
<connection>
<GID>433</GID>
<name>OUT_0</name></connection>
<connection>
<GID>422</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>826 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-155,-63.5,-155</points>
<connection>
<GID>593</GID>
<name>IN_0</name></connection>
<intersection>-63.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-63.5,-155,-63.5,-155</points>
<connection>
<GID>508</GID>
<name>IN_0</name></connection>
<intersection>-155 1</intersection></vsegment></shape></wire>
<wire>
<ID>673 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-75,93,-75</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<connection>
<GID>384</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>674 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-77,93,-77</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<intersection>93 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>93,-77,93,-77</points>
<connection>
<GID>384</GID>
<name>IN_1</name></connection>
<intersection>-77 1</intersection></vsegment></shape></wire>
<wire>
<ID>675 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-80,93,-80</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<connection>
<GID>416</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>676 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-82,93,-82</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<connection>
<GID>416</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>678 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-57,93,-57</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<intersection>93 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>93,-57,93,-57</points>
<connection>
<GID>383</GID>
<name>IN_1</name></connection>
<intersection>-57 1</intersection></vsegment></shape></wire>
<wire>
<ID>824 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-150,-53,-150</points>
<connection>
<GID>592</GID>
<name>IN_0</name></connection>
<intersection>-53 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-53,-150,-53,-150</points>
<connection>
<GID>587</GID>
<name>IN_1</name></connection>
<intersection>-150 1</intersection></vsegment></shape></wire>
<wire>
<ID>679 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157.5,-52,166,-52</points>
<connection>
<GID>443</GID>
<name>OUT</name></connection>
<connection>
<GID>442</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>680 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-50,157,-48</points>
<intersection>-50 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-50,166,-50</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-48,157,-48</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment></shape></wire>
<wire>
<ID>682 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-53,151.5,-53</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>151.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>151.5,-53,151.5,-53</points>
<connection>
<GID>443</GID>
<name>IN_1</name></connection>
<intersection>-53 1</intersection></vsegment></shape></wire>
<wire>
<ID>683 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-55,166,-55</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<connection>
<GID>440</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>684 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-81,185,-69</points>
<intersection>-81 2</intersection>
<intersection>-70 1</intersection>
<intersection>-69 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-70,194.5,-70</points>
<connection>
<GID>387</GID>
<name>IN_4</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-81,185,-81</points>
<connection>
<GID>439</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>185,-69,194.5,-69</points>
<connection>
<GID>387</GID>
<name>IN_5</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>686 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-71,183,-67</points>
<intersection>-71 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183,-67,194.5,-67</points>
<connection>
<GID>387</GID>
<name>IN_7</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-71,183,-71</points>
<connection>
<GID>447</GID>
<name>OUT</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>687 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-66,194.5,-66</points>
<connection>
<GID>446</GID>
<name>OUT</name></connection>
<connection>
<GID>387</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>688 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-65,183,-61</points>
<intersection>-65 1</intersection>
<intersection>-61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183,-65,194.5,-65</points>
<connection>
<GID>387</GID>
<name>IN_2</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-61,183,-61</points>
<connection>
<GID>444</GID>
<name>OUT</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>689 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-64,184,-56</points>
<intersection>-64 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172,-56,184,-56</points>
<connection>
<GID>440</GID>
<name>OUT</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184,-64,194.5,-64</points>
<connection>
<GID>387</GID>
<name>IN_1</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>690 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-63,185,-51</points>
<intersection>-63 1</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-63,194.5,-63</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-51,185,-51</points>
<connection>
<GID>442</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>691 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-62,166,-62</points>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>166 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>166,-62,166,-62</points>
<connection>
<GID>444</GID>
<name>IN_1</name></connection>
<intersection>-62 1</intersection></vsegment></shape></wire>
<wire>
<ID>692 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-60,166,-60</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<connection>
<GID>444</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>698 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-65,166,-65</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<connection>
<GID>446</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>699 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-67,166,-67</points>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<intersection>166 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>166,-67,166,-67</points>
<connection>
<GID>446</GID>
<name>IN_1</name></connection>
<intersection>-67 1</intersection></vsegment></shape></wire>
<wire>
<ID>700 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-70,166,-70</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<connection>
<GID>447</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>701 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>151,-72,155.5,-72</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>155.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>155.5,-72,155.5,-72</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<intersection>-72 3</intersection></vsegment></shape></wire>
<wire>
<ID>702 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>159.5,-72,166,-72</points>
<connection>
<GID>457</GID>
<name>OUT_0</name></connection>
<connection>
<GID>447</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>703 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-75,166,-75</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<connection>
<GID>448</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>704 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-77,166,-77</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>166 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>166,-77,166,-77</points>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<intersection>-77 1</intersection></vsegment></shape></wire>
<wire>
<ID>858 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-140,20,-140</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-140,20,-140</points>
<connection>
<GID>603</GID>
<name>IN_1</name></connection>
<intersection>-140 1</intersection></vsegment></shape></wire>
<wire>
<ID>705 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-80,166,-80</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<connection>
<GID>439</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>706 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-82,166,-82</points>
<connection>
<GID>439</GID>
<name>IN_1</name></connection>
<connection>
<GID>388</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>868 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-148,110,-144</points>
<intersection>-148 1</intersection>
<intersection>-144 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-148,121.5,-148</points>
<connection>
<GID>634</GID>
<name>IN_2</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-144,110,-144</points>
<connection>
<GID>582</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>707 </ID>
<shape>
<hsegment>
<ID>11</ID>
<points>201.5,-66.5,203.5,-66.5</points>
<connection>
<GID>460</GID>
<name>IN_0</name></connection>
<intersection>201.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>201.5,-66.5,201.5,-66.5</points>
<connection>
<GID>387</GID>
<name>OUT</name></connection>
<intersection>-66.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>862 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-136,78.5,-136</points>
<connection>
<GID>632</GID>
<name>IN_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-136,78.5,-136</points>
<connection>
<GID>627</GID>
<name>IN_1</name></connection>
<intersection>-136 1</intersection></vsegment></shape></wire>
<wire>
<ID>709 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-61.5,-94,-53,-94</points>
<connection>
<GID>466</GID>
<name>OUT</name></connection>
<connection>
<GID>465</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>710 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-92,-62,-90</points>
<intersection>-92 1</intersection>
<intersection>-90 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-92,-53,-92</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-68,-90,-62,-90</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>856 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-165,20,-165</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<connection>
<GID>602</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>711 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-93,-67.5,-93</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<intersection>-67.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-67.5,-93,-67.5,-93</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>866 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-154,110,-150</points>
<intersection>-154 2</intersection>
<intersection>-150 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-150,121.5,-150</points>
<connection>
<GID>634</GID>
<name>IN_7</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-154,110,-154</points>
<connection>
<GID>630</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>713 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-97,-53,-97</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<connection>
<GID>463</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>714 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-123,-34,-111</points>
<intersection>-123 2</intersection>
<intersection>-112 1</intersection>
<intersection>-111 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-112,-24.5,-112</points>
<connection>
<GID>477</GID>
<name>IN_4</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-123,-34,-123</points>
<connection>
<GID>462</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-34,-111,-24.5,-111</points>
<connection>
<GID>477</GID>
<name>IN_5</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>876 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>78,-155,82.5,-155</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>82.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>82.5,-155,82.5,-155</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>-155 3</intersection></vsegment></shape></wire>
<wire>
<ID>715 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-118,-35,-110</points>
<intersection>-118 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,-110,-24.5,-110</points>
<connection>
<GID>477</GID>
<name>IN_6</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-118,-35,-118</points>
<connection>
<GID>472</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>870 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-146,112,-134</points>
<intersection>-146 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-146,121.5,-146</points>
<connection>
<GID>634</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-134,112,-134</points>
<connection>
<GID>626</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>717 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-108,-24.5,-108</points>
<connection>
<GID>469</GID>
<name>OUT</name></connection>
<connection>
<GID>477</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>718 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-107,-36,-103</points>
<intersection>-107 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-107,-24.5,-107</points>
<connection>
<GID>477</GID>
<name>IN_2</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-103,-36,-103</points>
<connection>
<GID>467</GID>
<name>OUT</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>864 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-164,112,-152</points>
<intersection>-164 2</intersection>
<intersection>-153 1</intersection>
<intersection>-152 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-153,121.5,-153</points>
<connection>
<GID>634</GID>
<name>IN_4</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-164,112,-164</points>
<connection>
<GID>624</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>112,-152,121.5,-152</points>
<connection>
<GID>634</GID>
<name>IN_5</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>719 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-106,-35,-98</points>
<intersection>-106 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-98,-35,-98</points>
<connection>
<GID>463</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-35,-106,-24.5,-106</points>
<connection>
<GID>477</GID>
<name>IN_1</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>720 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-105,-34,-93</points>
<intersection>-105 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-105,-24.5,-105</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-93,-34,-93</points>
<connection>
<GID>465</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>874 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-150,93,-150</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-150,93,-150</points>
<connection>
<GID>629</GID>
<name>IN_1</name></connection>
<intersection>-150 1</intersection></vsegment></shape></wire>
<wire>
<ID>721 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-104,-53,-104</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>-53 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-53,-104,-53,-104</points>
<connection>
<GID>467</GID>
<name>IN_1</name></connection>
<intersection>-104 1</intersection></vsegment></shape></wire>
<wire>
<ID>722 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-102,-53,-102</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<connection>
<GID>467</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>724 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-109,-53,-109</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>-53 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-53,-109,-53,-109</points>
<connection>
<GID>469</GID>
<name>IN_1</name></connection>
<intersection>-109 1</intersection></vsegment></shape></wire>
<wire>
<ID>878 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-158,93,-158</points>
<connection>
<GID>642</GID>
<name>IN_0</name></connection>
<connection>
<GID>597</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>725 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-112,-53,-112</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<connection>
<GID>471</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>726 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-114,-63.5,-114</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>-63.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-63.5,-114,-63.5,-114</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>-114 1</intersection></vsegment></shape></wire>
<wire>
<ID>872 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-143,93,-143</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<connection>
<GID>582</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>727 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-114,-53,-114</points>
<connection>
<GID>487</GID>
<name>OUT_0</name></connection>
<connection>
<GID>471</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>882 </ID>
<shape>
<hsegment>
<ID>11</ID>
<points>128.5,-149.5,130.5,-149.5</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>128.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>128.5,-149.5,128.5,-149.5</points>
<connection>
<GID>634</GID>
<name>OUT</name></connection>
<intersection>-149.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>729 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-119,-53,-119</points>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<intersection>-53 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-53,-119,-53,-119</points>
<connection>
<GID>472</GID>
<name>IN_1</name></connection>
<intersection>-119 1</intersection></vsegment></shape></wire>
<wire>
<ID>730 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-122,-53,-122</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<connection>
<GID>462</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>886 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-134,151.5,-134</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>151.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>151.5,-134,151.5,-134</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>-134 1</intersection></vsegment></shape></wire>
<wire>
<ID>733 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-99,-53,-99</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>-53 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-53,-99,-53,-99</points>
<connection>
<GID>463</GID>
<name>IN_1</name></connection>
<intersection>-99 1</intersection></vsegment></shape></wire>
<wire>
<ID>734 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-94,20,-94</points>
<connection>
<GID>515</GID>
<name>OUT</name></connection>
<connection>
<GID>513</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>880 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-163,93,-163</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<connection>
<GID>624</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>735 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-92,11,-90</points>
<intersection>-92 1</intersection>
<intersection>-90 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-92,20,-92</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-90,11,-90</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>890 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-159,184,-151</points>
<intersection>-159 2</intersection>
<intersection>-151 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-151,194.5,-151</points>
<connection>
<GID>599</GID>
<name>IN_6</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-159,184,-159</points>
<connection>
<GID>656</GID>
<name>OUT</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>737 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-95,5.5,-95</points>
<connection>
<GID>522</GID>
<name>IN_0</name></connection>
<intersection>5.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5.5,-95,5.5,-95</points>
<connection>
<GID>515</GID>
<name>IN_1</name></connection>
<intersection>-95 1</intersection></vsegment></shape></wire>
<wire>
<ID>738 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-97,20,-97</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<connection>
<GID>510</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>894 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-147,184,-139</points>
<intersection>-147 2</intersection>
<intersection>-139 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172,-139,184,-139</points>
<connection>
<GID>648</GID>
<name>OUT</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184,-147,194.5,-147</points>
<connection>
<GID>599</GID>
<name>IN_1</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>741 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-113,37,-109</points>
<intersection>-113 2</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-109,48.5,-109</points>
<connection>
<GID>524</GID>
<name>IN_7</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-113,37,-113</points>
<connection>
<GID>519</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>742 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-108,48.5,-108</points>
<connection>
<GID>518</GID>
<name>OUT</name></connection>
<connection>
<GID>524</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>744 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-106,38,-98</points>
<intersection>-106 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-98,38,-98</points>
<connection>
<GID>510</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-106,48.5,-106</points>
<connection>
<GID>524</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>770 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-105,112,-93</points>
<intersection>-105 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-105,121.5,-105</points>
<connection>
<GID>547</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-93,112,-93</points>
<connection>
<GID>539</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>745 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-105,39,-93</points>
<intersection>-105 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-105,48.5,-105</points>
<connection>
<GID>524</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-93,39,-93</points>
<connection>
<GID>513</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>746 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-104,20,-104</points>
<connection>
<GID>526</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-104,20,-104</points>
<connection>
<GID>516</GID>
<name>IN_1</name></connection>
<intersection>-104 1</intersection></vsegment></shape></wire>
<wire>
<ID>780 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-122,93,-122</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<connection>
<GID>537</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>747 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-102,20,-102</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<connection>
<GID>516</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>774 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-109,93,-109</points>
<connection>
<GID>551</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-109,93,-109</points>
<connection>
<GID>542</GID>
<name>IN_1</name></connection>
<intersection>-109 1</intersection></vsegment></shape></wire>
<wire>
<ID>749 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-109,20,-109</points>
<connection>
<GID>528</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-109,20,-109</points>
<connection>
<GID>518</GID>
<name>IN_1</name></connection>
<intersection>-109 1</intersection></vsegment></shape></wire>
<wire>
<ID>750 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-112,20,-112</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<connection>
<GID>519</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>778 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-117,93,-117</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<connection>
<GID>493</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>753 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-117,20,-117</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<connection>
<GID>520</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>754 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-119,20,-119</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-119,20,-119</points>
<connection>
<GID>520</GID>
<name>IN_1</name></connection>
<intersection>-119 1</intersection></vsegment></shape></wire>
<wire>
<ID>788 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-97,166,-97</points>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<connection>
<GID>561</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>755 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-122,20,-122</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<connection>
<GID>509</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>756 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-124,20,-124</points>
<connection>
<GID>534</GID>
<name>IN_0</name></connection>
<connection>
<GID>509</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>782 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>128.5,-108.5,130.5,-108.5</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<intersection>128.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>128.5,-108.5,128.5,-108.5</points>
<connection>
<GID>547</GID>
<name>OUT</name></connection>
<intersection>-108.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>757 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-108.5,57.5,-108.5</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>55.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>55.5,-108.5,55.5,-108.5</points>
<connection>
<GID>524</GID>
<name>OUT</name></connection>
<intersection>-108.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>758 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-99,20,-99</points>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-99,20,-99</points>
<connection>
<GID>510</GID>
<name>IN_1</name></connection>
<intersection>-99 1</intersection></vsegment></shape></wire>
<wire>
<ID>760 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-92,84,-90</points>
<intersection>-92 1</intersection>
<intersection>-90 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-92,93,-92</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-90,84,-90</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>786 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-93,151.5,-93</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<intersection>151.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>151.5,-93,151.5,-93</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>761 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-93,78.5,-93</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-93,78.5,-93</points>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>762 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-95,78.5,-95</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-95,78.5,-95</points>
<connection>
<GID>540</GID>
<name>IN_1</name></connection>
<intersection>-95 1</intersection></vsegment></shape></wire>
<wire>
<ID>796 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-104,166,-104</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-104,166,-104</points>
<connection>
<GID>565</GID>
<name>IN_1</name></connection>
<intersection>-104 1</intersection></vsegment></shape></wire>
<wire>
<ID>763 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-97,93,-97</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<connection>
<GID>492</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>764 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-123,112,-111</points>
<intersection>-123 2</intersection>
<intersection>-112 1</intersection>
<intersection>-111 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-112,121.5,-112</points>
<connection>
<GID>547</GID>
<name>IN_4</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-123,112,-123</points>
<connection>
<GID>537</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>112,-111,121.5,-111</points>
<connection>
<GID>547</GID>
<name>IN_5</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>790 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-118,184,-110</points>
<intersection>-118 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-110,194.5,-110</points>
<connection>
<GID>496</GID>
<name>IN_6</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-118,184,-118</points>
<connection>
<GID>569</GID>
<name>OUT</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>765 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-118,111,-110</points>
<intersection>-118 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-110,121.5,-110</points>
<connection>
<GID>547</GID>
<name>IN_6</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-118,111,-118</points>
<connection>
<GID>493</GID>
<name>OUT</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>766 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-113,110,-109</points>
<intersection>-113 2</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-109,121.5,-109</points>
<connection>
<GID>547</GID>
<name>IN_7</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-113,110,-113</points>
<connection>
<GID>543</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>784 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157.5,-94,166,-94</points>
<connection>
<GID>564</GID>
<name>OUT</name></connection>
<connection>
<GID>563</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>767 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99,-108,121.5,-108</points>
<connection>
<GID>542</GID>
<name>OUT</name></connection>
<connection>
<GID>547</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>785 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-92,157,-90</points>
<intersection>-92 1</intersection>
<intersection>-90 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-92,166,-92</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-90,157,-90</points>
<connection>
<GID>566</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment></shape></wire>
<wire>
<ID>787 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-95,151.5,-95</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>151.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>151.5,-95,151.5,-95</points>
<connection>
<GID>564</GID>
<name>IN_1</name></connection>
<intersection>-95 1</intersection></vsegment></shape></wire>
<wire>
<ID>789 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-123,185,-111</points>
<intersection>-123 2</intersection>
<intersection>-112 1</intersection>
<intersection>-111 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-112,194.5,-112</points>
<connection>
<GID>496</GID>
<name>IN_4</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-123,185,-123</points>
<connection>
<GID>560</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>185,-111,194.5,-111</points>
<connection>
<GID>496</GID>
<name>IN_5</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>793 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-107,183,-103</points>
<intersection>-107 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183,-107,194.5,-107</points>
<connection>
<GID>496</GID>
<name>IN_2</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-103,183,-103</points>
<connection>
<GID>565</GID>
<name>OUT</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>797 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-102,166,-102</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<connection>
<GID>565</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>801 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>151,-114,155.5,-114</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>155.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>155.5,-114,155.5,-114</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<intersection>-114 3</intersection></vsegment></shape></wire>
<wire>
<ID>805 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-122,166,-122</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<connection>
<GID>560</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>808 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-99,166,-99</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-99,166,-99</points>
<connection>
<GID>561</GID>
<name>IN_1</name></connection>
<intersection>-99 1</intersection></vsegment></shape></wire>
<wire>
<ID>809 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-61.5,-135,-53,-135</points>
<connection>
<GID>585</GID>
<name>OUT</name></connection>
<connection>
<GID>584</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>810 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-133,-62,-131</points>
<intersection>-133 1</intersection>
<intersection>-131 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-133,-53,-133</points>
<connection>
<GID>584</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-68,-131,-62,-131</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>811 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-68,-134,-67.5,-134</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>-67.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-67.5,-134,-67.5,-134</points>
<connection>
<GID>585</GID>
<name>IN_0</name></connection>
<intersection>-134 3</intersection></vsegment></shape></wire>
<wire>
<ID>813 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-138,-53,-138</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<connection>
<GID>583</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>814 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-164,-34,-152</points>
<intersection>-164 2</intersection>
<intersection>-153 1</intersection>
<intersection>-152 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-153,-24.5,-153</points>
<connection>
<GID>590</GID>
<name>IN_4</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-164,-34,-164</points>
<connection>
<GID>499</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-34,-152,-24.5,-152</points>
<connection>
<GID>590</GID>
<name>IN_5</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>817 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-149,-24.5,-149</points>
<connection>
<GID>587</GID>
<name>OUT</name></connection>
<connection>
<GID>590</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>818 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-148,-36,-144</points>
<intersection>-148 1</intersection>
<intersection>-144 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-148,-24.5,-148</points>
<connection>
<GID>590</GID>
<name>IN_2</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-144,-36,-144</points>
<connection>
<GID>586</GID>
<name>OUT</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>819 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-147,-35,-139</points>
<intersection>-147 2</intersection>
<intersection>-139 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-139,-35,-139</points>
<connection>
<GID>583</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-35,-147,-24.5,-147</points>
<connection>
<GID>590</GID>
<name>IN_1</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>820 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-146,-34,-134</points>
<intersection>-146 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-146,-24.5,-146</points>
<connection>
<GID>590</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-134,-34,-134</points>
<connection>
<GID>584</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>821 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-145,-53,-145</points>
<connection>
<GID>591</GID>
<name>IN_0</name></connection>
<intersection>-53 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-53,-145,-53,-145</points>
<connection>
<GID>586</GID>
<name>IN_1</name></connection>
<intersection>-145 1</intersection></vsegment></shape></wire>
<wire>
<ID>823 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-148,-53,-148</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<connection>
<GID>587</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>827 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-155,-53,-155</points>
<connection>
<GID>508</GID>
<name>OUT_0</name></connection>
<connection>
<GID>502</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>828 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-158,-53,-158</points>
<connection>
<GID>594</GID>
<name>IN_0</name></connection>
<connection>
<GID>588</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>829 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-160,-53,-160</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<intersection>-53 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-53,-160,-53,-160</points>
<connection>
<GID>588</GID>
<name>IN_1</name></connection>
<intersection>-160 1</intersection></vsegment></shape></wire>
<wire>
<ID>831 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-165,-53,-165</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<connection>
<GID>499</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>832 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-149.5,-15.5,-149.5</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>-17.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-17.5,-149.5,-17.5,-149.5</points>
<connection>
<GID>590</GID>
<name>OUT</name></connection>
<intersection>-149.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>833 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-140,-53,-140</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<intersection>-53 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-53,-140,-53,-140</points>
<connection>
<GID>583</GID>
<name>IN_1</name></connection>
<intersection>-140 1</intersection></vsegment></shape></wire>
<wire>
<ID>834 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-135,20,-135</points>
<connection>
<GID>606</GID>
<name>OUT</name></connection>
<connection>
<GID>605</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>835 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-133,11,-131</points>
<intersection>-133 1</intersection>
<intersection>-131 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-133,20,-133</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-131,11,-131</points>
<connection>
<GID>608</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>836 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-134,5.5,-134</points>
<connection>
<GID>611</GID>
<name>IN_0</name></connection>
<intersection>5.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5.5,-134,5.5,-134</points>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<intersection>-134 1</intersection></vsegment></shape></wire>
<wire>
<ID>837 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-136,5.5,-136</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>5.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5.5,-136,5.5,-136</points>
<connection>
<GID>606</GID>
<name>IN_1</name></connection>
<intersection>-136 1</intersection></vsegment></shape></wire>
<wire>
<ID>838 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-138,20,-138</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<connection>
<GID>603</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>839 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-164,39,-152</points>
<intersection>-164 2</intersection>
<intersection>-153 1</intersection>
<intersection>-152 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-153,48.5,-153</points>
<connection>
<GID>614</GID>
<name>IN_4</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-164,39,-164</points>
<connection>
<GID>602</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>39,-152,48.5,-152</points>
<connection>
<GID>614</GID>
<name>IN_5</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>840 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-159,38,-151</points>
<intersection>-159 2</intersection>
<intersection>-151 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-151,48.5,-151</points>
<connection>
<GID>614</GID>
<name>IN_6</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-159,38,-159</points>
<connection>
<GID>610</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>841 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-154,37,-150</points>
<intersection>-154 2</intersection>
<intersection>-150 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-150,48.5,-150</points>
<connection>
<GID>614</GID>
<name>IN_7</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-154,37,-154</points>
<connection>
<GID>609</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>842 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-149,48.5,-149</points>
<connection>
<GID>474</GID>
<name>OUT</name></connection>
<connection>
<GID>614</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>843 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-148,37,-144</points>
<intersection>-148 1</intersection>
<intersection>-144 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-148,48.5,-148</points>
<connection>
<GID>614</GID>
<name>IN_2</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-144,37,-144</points>
<connection>
<GID>607</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>844 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-147,38,-139</points>
<intersection>-147 2</intersection>
<intersection>-139 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-139,38,-139</points>
<connection>
<GID>603</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-147,48.5,-147</points>
<connection>
<GID>614</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>845 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-146,39,-134</points>
<intersection>-146 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-146,48.5,-146</points>
<connection>
<GID>614</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-134,39,-134</points>
<connection>
<GID>605</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>846 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-145,20,-145</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-145,20,-145</points>
<connection>
<GID>607</GID>
<name>IN_1</name></connection>
<intersection>-145 1</intersection></vsegment></shape></wire>
<wire>
<ID>847 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-143,20,-143</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<connection>
<GID>607</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>849 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-150,20,-150</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-150,20,-150</points>
<connection>
<GID>474</GID>
<name>IN_1</name></connection>
<intersection>-150 1</intersection></vsegment></shape></wire>
<wire>
<ID>850 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-153,20,-153</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<connection>
<GID>609</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>851 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-155,9.5,-155</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<intersection>9.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>9.5,-155,9.5,-155</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<intersection>-155 1</intersection></vsegment></shape></wire>
<wire>
<ID>852 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-155,20,-155</points>
<connection>
<GID>619</GID>
<name>OUT_0</name></connection>
<connection>
<GID>609</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>853 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-158,20,-158</points>
<connection>
<GID>620</GID>
<name>IN_0</name></connection>
<connection>
<GID>610</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>854 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-160,20,-160</points>
<connection>
<GID>621</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-160,20,-160</points>
<connection>
<GID>610</GID>
<name>IN_1</name></connection>
<intersection>-160 1</intersection></vsegment></shape></wire>
<wire>
<ID>855 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-163,20,-163</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<connection>
<GID>602</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>857 </ID>
<shape>
<hsegment>
<ID>9</ID>
<points>55.5,-149.5,57.5,-149.5</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<intersection>55.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>55.5,-149.5,55.5,-149.5</points>
<connection>
<GID>614</GID>
<name>OUT</name></connection>
<intersection>-149.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>859 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-135,93,-135</points>
<connection>
<GID>627</GID>
<name>OUT</name></connection>
<connection>
<GID>626</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>860 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-133,84,-131</points>
<intersection>-133 1</intersection>
<intersection>-131 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-133,93,-133</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-131,84,-131</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>861 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-134,78.5,-134</points>
<connection>
<GID>631</GID>
<name>IN_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-134,78.5,-134</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>-134 1</intersection></vsegment></shape></wire>
<wire>
<ID>863 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-138,93,-138</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<connection>
<GID>596</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>865 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-159,111,-151</points>
<intersection>-159 2</intersection>
<intersection>-151 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-151,121.5,-151</points>
<connection>
<GID>634</GID>
<name>IN_6</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-159,111,-159</points>
<connection>
<GID>597</GID>
<name>OUT</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>867 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99,-149,121.5,-149</points>
<connection>
<GID>629</GID>
<name>OUT</name></connection>
<connection>
<GID>634</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>869 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-147,111,-139</points>
<intersection>-147 2</intersection>
<intersection>-139 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-139,111,-139</points>
<connection>
<GID>596</GID>
<name>OUT</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111,-147,121.5,-147</points>
<connection>
<GID>634</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>871 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-145,93,-145</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-145,93,-145</points>
<connection>
<GID>582</GID>
<name>IN_1</name></connection>
<intersection>-145 1</intersection></vsegment></shape></wire>
<wire>
<ID>873 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-148,93,-148</points>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<connection>
<GID>629</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>875 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-153,93,-153</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<connection>
<GID>630</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>877 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-155,93,-155</points>
<connection>
<GID>641</GID>
<name>OUT_0</name></connection>
<connection>
<GID>630</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>879 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-160,93,-160</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-160,93,-160</points>
<connection>
<GID>597</GID>
<name>IN_1</name></connection>
<intersection>-160 1</intersection></vsegment></shape></wire>
<wire>
<ID>887 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-136,151.5,-136</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>151.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>151.5,-136,151.5,-136</points>
<connection>
<GID>651</GID>
<name>IN_1</name></connection>
<intersection>-136 1</intersection></vsegment></shape></wire>
<wire>
<ID>895 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-146,185,-134</points>
<intersection>-146 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-146,194.5,-146</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-134,185,-134</points>
<connection>
<GID>650</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>896 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-145,166,-145</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-145,166,-145</points>
<connection>
<GID>652</GID>
<name>IN_1</name></connection>
<intersection>-145 1</intersection></vsegment></shape></wire>
<wire>
<ID>900 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-153,166,-153</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<connection>
<GID>655</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>902 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>159.5,-155,166,-155</points>
<connection>
<GID>665</GID>
<name>OUT_0</name></connection>
<connection>
<GID>655</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>904 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-160,166,-160</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-160,166,-160</points>
<connection>
<GID>656</GID>
<name>IN_1</name></connection>
<intersection>-160 1</intersection></vsegment></shape></wire>
<wire>
<ID>907 </ID>
<shape>
<hsegment>
<ID>11</ID>
<points>201.5,-149.5,203.5,-149.5</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>201.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>201.5,-149.5,201.5,-149.5</points>
<connection>
<GID>599</GID>
<name>OUT</name></connection>
<intersection>-149.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>908 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-140,166,-140</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-140,166,-140</points>
<connection>
<GID>648</GID>
<name>IN_1</name></connection>
<intersection>-140 1</intersection></vsegment></shape></wire></page 1></circuit>