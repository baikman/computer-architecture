
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-32.95,39.6893,61.95,-63.2229</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>14.5,-13</position>
<gparam>LABEL_TEXT Go to https://cedar.to/vjyQw7 to download the latest version!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>14.5,-9.5</position>
<gparam>LABEL_TEXT Error: This file was made with a newer version of Cedar Logic!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 0>
</circuit>
<throw_away></throw_away>

	<version>2.3.5 | 2018-09-25 23:06:05</version><circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-106.394,0.149845,101.131,-104.545</PageViewport>
<gate>
<ID>2</ID>
<type>AI_RAM_12x16</type>
<position>23,12.5</position>
<input>
<ID>ADDRESS_0</ID>197 </input>
<input>
<ID>ADDRESS_1</ID>198 </input>
<input>
<ID>ADDRESS_10</ID>203 </input>
<input>
<ID>ADDRESS_11</ID>204 </input>
<input>
<ID>ADDRESS_2</ID>195 </input>
<input>
<ID>ADDRESS_3</ID>201 </input>
<input>
<ID>ADDRESS_4</ID>199 </input>
<input>
<ID>ADDRESS_5</ID>202 </input>
<input>
<ID>ADDRESS_6</ID>200 </input>
<input>
<ID>ADDRESS_7</ID>193 </input>
<input>
<ID>ADDRESS_8</ID>194 </input>
<input>
<ID>ADDRESS_9</ID>196 </input>
<input>
<ID>DATA_IN_0</ID>6 </input>
<input>
<ID>DATA_IN_1</ID>7 </input>
<input>
<ID>DATA_IN_10</ID>13 </input>
<input>
<ID>DATA_IN_11</ID>15 </input>
<input>
<ID>DATA_IN_12</ID>10 </input>
<input>
<ID>DATA_IN_13</ID>9 </input>
<input>
<ID>DATA_IN_14</ID>12 </input>
<input>
<ID>DATA_IN_15</ID>17 </input>
<input>
<ID>DATA_IN_2</ID>2 </input>
<input>
<ID>DATA_IN_3</ID>3 </input>
<input>
<ID>DATA_IN_4</ID>4 </input>
<input>
<ID>DATA_IN_5</ID>8 </input>
<input>
<ID>DATA_IN_6</ID>5 </input>
<input>
<ID>DATA_IN_7</ID>11 </input>
<input>
<ID>DATA_IN_8</ID>16 </input>
<input>
<ID>DATA_IN_9</ID>14 </input>
<output>
<ID>DATA_OUT_0</ID>6 </output>
<output>
<ID>DATA_OUT_1</ID>7 </output>
<output>
<ID>DATA_OUT_10</ID>13 </output>
<output>
<ID>DATA_OUT_11</ID>15 </output>
<output>
<ID>DATA_OUT_12</ID>10 </output>
<output>
<ID>DATA_OUT_13</ID>9 </output>
<output>
<ID>DATA_OUT_14</ID>12 </output>
<output>
<ID>DATA_OUT_15</ID>17 </output>
<output>
<ID>DATA_OUT_2</ID>2 </output>
<output>
<ID>DATA_OUT_3</ID>3 </output>
<output>
<ID>DATA_OUT_4</ID>4 </output>
<output>
<ID>DATA_OUT_5</ID>8 </output>
<output>
<ID>DATA_OUT_6</ID>5 </output>
<output>
<ID>DATA_OUT_7</ID>11 </output>
<output>
<ID>DATA_OUT_8</ID>16 </output>
<output>
<ID>DATA_OUT_9</ID>14 </output>
<input>
<ID>ENABLE_0</ID>564 </input>
<input>
<ID>write_clock</ID>491 </input>
<input>
<ID>write_enable</ID>563 </input>
<gparam>angle 0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>34.5,14</position>
<input>
<ID>IN_0</ID>491 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>0,-17.5</position>
<gparam>LABEL_TEXT Address Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AE_REGISTER8</type>
<position>3.5,-148.5</position>
<input>
<ID>IN_0</ID>609 </input>
<input>
<ID>IN_1</ID>610 </input>
<input>
<ID>IN_2</ID>611 </input>
<input>
<ID>IN_3</ID>614 </input>
<input>
<ID>IN_4</ID>615 </input>
<input>
<ID>IN_5</ID>616 </input>
<input>
<ID>IN_6</ID>612 </input>
<input>
<ID>IN_7</ID>613 </input>
<input>
<ID>clock</ID>493 </input>
<input>
<ID>count_up</ID>581 </input>
<input>
<ID>load</ID>591 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>76</ID>
<type>DE_TO</type>
<position>-7,4.5</position>
<input>
<ID>IN_0</ID>492 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>12</ID>
<type>AI_REGISTER12</type>
<position>40,-53</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>107 </input>
<input>
<ID>IN_10</ID>106 </input>
<input>
<ID>IN_11</ID>101 </input>
<input>
<ID>IN_2</ID>109 </input>
<input>
<ID>IN_3</ID>110 </input>
<input>
<ID>IN_4</ID>99 </input>
<input>
<ID>IN_5</ID>104 </input>
<input>
<ID>IN_6</ID>105 </input>
<input>
<ID>IN_7</ID>100 </input>
<input>
<ID>IN_8</ID>103 </input>
<input>
<ID>IN_9</ID>102 </input>
<output>
<ID>OUT_0</ID>552 </output>
<output>
<ID>OUT_1</ID>557 </output>
<output>
<ID>OUT_10</ID>561 </output>
<output>
<ID>OUT_11</ID>562 </output>
<output>
<ID>OUT_2</ID>551 </output>
<output>
<ID>OUT_3</ID>556 </output>
<output>
<ID>OUT_4</ID>553 </output>
<output>
<ID>OUT_5</ID>554 </output>
<output>
<ID>OUT_6</ID>555 </output>
<output>
<ID>OUT_7</ID>558 </output>
<output>
<ID>OUT_8</ID>559 </output>
<output>
<ID>OUT_9</ID>560 </output>
<input>
<ID>clear</ID>569 </input>
<input>
<ID>clock</ID>498 </input>
<input>
<ID>count_enable</ID>572 </input>
<input>
<ID>count_up</ID>571 </input>
<input>
<ID>load</ID>570 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>14</ID>
<type>AM_REGISTER16</type>
<position>36,-90</position>
<input>
<ID>IN_0</ID>254 </input>
<input>
<ID>IN_1</ID>255 </input>
<input>
<ID>IN_10</ID>261 </input>
<input>
<ID>IN_11</ID>266 </input>
<input>
<ID>IN_12</ID>262 </input>
<input>
<ID>IN_13</ID>265 </input>
<input>
<ID>IN_14</ID>263 </input>
<input>
<ID>IN_15</ID>264 </input>
<input>
<ID>IN_2</ID>256 </input>
<input>
<ID>IN_3</ID>257 </input>
<input>
<ID>IN_4</ID>258 </input>
<input>
<ID>IN_5</ID>269 </input>
<input>
<ID>IN_6</ID>259 </input>
<input>
<ID>IN_7</ID>268 </input>
<input>
<ID>IN_8</ID>260 </input>
<input>
<ID>IN_9</ID>267 </input>
<output>
<ID>OUT_0</ID>414 </output>
<output>
<ID>OUT_1</ID>399 </output>
<output>
<ID>OUT_10</ID>405 </output>
<output>
<ID>OUT_11</ID>403 </output>
<output>
<ID>OUT_12</ID>404 </output>
<output>
<ID>OUT_13</ID>406 </output>
<output>
<ID>OUT_14</ID>407 </output>
<output>
<ID>OUT_15</ID>409 </output>
<output>
<ID>OUT_2</ID>410 </output>
<output>
<ID>OUT_3</ID>400 </output>
<output>
<ID>OUT_4</ID>401 </output>
<output>
<ID>OUT_5</ID>408 </output>
<output>
<ID>OUT_6</ID>411 </output>
<output>
<ID>OUT_7</ID>412 </output>
<output>
<ID>OUT_8</ID>402 </output>
<output>
<ID>OUT_9</ID>413 </output>
<input>
<ID>clear</ID>583 </input>
<input>
<ID>clock</ID>496 </input>
<input>
<ID>count_enable</ID>577 </input>
<input>
<ID>count_up</ID>578 </input>
<input>
<ID>load</ID>582 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>-1,-158</position>
<input>
<ID>IN_0</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>6</ID>
<type>AI_REGISTER12</type>
<position>-1,-31.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>179 </input>
<input>
<ID>IN_10</ID>177 </input>
<input>
<ID>IN_11</ID>178 </input>
<input>
<ID>IN_2</ID>93 </input>
<input>
<ID>IN_3</ID>96 </input>
<input>
<ID>IN_4</ID>97 </input>
<input>
<ID>IN_5</ID>98 </input>
<input>
<ID>IN_6</ID>176 </input>
<input>
<ID>IN_7</ID>94 </input>
<input>
<ID>IN_8</ID>180 </input>
<input>
<ID>IN_9</ID>175 </input>
<output>
<ID>OUT_0</ID>188 </output>
<output>
<ID>OUT_1</ID>182 </output>
<output>
<ID>OUT_10</ID>191 </output>
<output>
<ID>OUT_11</ID>192 </output>
<output>
<ID>OUT_2</ID>190 </output>
<output>
<ID>OUT_3</ID>189 </output>
<output>
<ID>OUT_4</ID>181 </output>
<output>
<ID>OUT_5</ID>183 </output>
<output>
<ID>OUT_6</ID>184 </output>
<output>
<ID>OUT_7</ID>185 </output>
<output>
<ID>OUT_8</ID>187 </output>
<output>
<ID>OUT_9</ID>186 </output>
<input>
<ID>clear</ID>565 </input>
<input>
<ID>clock</ID>499 </input>
<input>
<ID>count_enable</ID>568 </input>
<input>
<ID>load</ID>566 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>8</ID>
<type>AM_REGISTER16</type>
<position>-6,-70.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>116 </input>
<input>
<ID>IN_10</ID>115 </input>
<input>
<ID>IN_11</ID>120 </input>
<input>
<ID>IN_12</ID>122 </input>
<input>
<ID>IN_13</ID>117 </input>
<input>
<ID>IN_14</ID>118 </input>
<input>
<ID>IN_15</ID>121 </input>
<input>
<ID>IN_2</ID>123 </input>
<input>
<ID>IN_3</ID>112 </input>
<input>
<ID>IN_4</ID>126 </input>
<input>
<ID>IN_5</ID>119 </input>
<input>
<ID>IN_6</ID>114 </input>
<input>
<ID>IN_7</ID>113 </input>
<input>
<ID>IN_8</ID>111 </input>
<input>
<ID>IN_9</ID>124 </input>
<output>
<ID>OUT_0</ID>369 </output>
<output>
<ID>OUT_1</ID>374 </output>
<output>
<ID>OUT_10</ID>377 </output>
<output>
<ID>OUT_11</ID>379 </output>
<output>
<ID>OUT_12</ID>380 </output>
<output>
<ID>OUT_13</ID>381 </output>
<output>
<ID>OUT_14</ID>371 </output>
<output>
<ID>OUT_15</ID>382 </output>
<output>
<ID>OUT_2</ID>375 </output>
<output>
<ID>OUT_3</ID>367 </output>
<output>
<ID>OUT_4</ID>373 </output>
<output>
<ID>OUT_5</ID>372 </output>
<output>
<ID>OUT_6</ID>368 </output>
<output>
<ID>OUT_7</ID>378 </output>
<output>
<ID>OUT_8</ID>370 </output>
<output>
<ID>OUT_9</ID>376 </output>
<input>
<ID>clear</ID>573 </input>
<input>
<ID>clock</ID>497 </input>
<input>
<ID>count_enable</ID>575 </input>
<input>
<ID>count_up</ID>574 </input>
<input>
<ID>load</ID>576 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>32.5,-39.5</position>
<gparam>LABEL_TEXT Program Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>-5.5,-54</position>
<gparam>LABEL_TEXT Data Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>36.5,-73.5</position>
<gparam>LABEL_TEXT Accumulator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>31.5,-144.5</position>
<input>
<ID>IN_0</ID>494 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>16</ID>
<type>AM_REGISTER16</type>
<position>-6.5,-111.5</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_10</ID>147 </input>
<input>
<ID>IN_11</ID>145 </input>
<input>
<ID>IN_12</ID>152 </input>
<input>
<ID>IN_13</ID>153 </input>
<input>
<ID>IN_14</ID>155 </input>
<input>
<ID>IN_15</ID>158 </input>
<input>
<ID>IN_2</ID>150 </input>
<input>
<ID>IN_3</ID>149 </input>
<input>
<ID>IN_4</ID>148 </input>
<input>
<ID>IN_5</ID>156 </input>
<input>
<ID>IN_6</ID>143 </input>
<input>
<ID>IN_7</ID>154 </input>
<input>
<ID>IN_8</ID>151 </input>
<input>
<ID>IN_9</ID>157 </input>
<output>
<ID>OUT_0</ID>431 </output>
<output>
<ID>OUT_1</ID>432 </output>
<output>
<ID>OUT_10</ID>439 </output>
<output>
<ID>OUT_11</ID>444 </output>
<output>
<ID>OUT_12</ID>443 </output>
<output>
<ID>OUT_13</ID>445 </output>
<output>
<ID>OUT_14</ID>442 </output>
<output>
<ID>OUT_15</ID>446 </output>
<output>
<ID>OUT_2</ID>433 </output>
<output>
<ID>OUT_3</ID>434 </output>
<output>
<ID>OUT_4</ID>435 </output>
<output>
<ID>OUT_5</ID>440 </output>
<output>
<ID>OUT_6</ID>441 </output>
<output>
<ID>OUT_7</ID>436 </output>
<output>
<ID>OUT_8</ID>437 </output>
<output>
<ID>OUT_9</ID>438 </output>
<input>
<ID>clock</ID>495 </input>
<input>
<ID>count_up</ID>579 </input>
<input>
<ID>load</ID>585 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>-10,-124.5</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>-6,-96.5</position>
<gparam>LABEL_TEXT Instruction Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>32,-102.5</position>
<input>
<ID>IN_0</ID>496 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>18</ID>
<type>AM_REGISTER16</type>
<position>35.5,-131.5</position>
<input>
<ID>IN_0</ID>164 </input>
<input>
<ID>IN_1</ID>168 </input>
<input>
<ID>IN_10</ID>171 </input>
<input>
<ID>IN_11</ID>172 </input>
<input>
<ID>IN_12</ID>174 </input>
<input>
<ID>IN_13</ID>159 </input>
<input>
<ID>IN_14</ID>162 </input>
<input>
<ID>IN_15</ID>163 </input>
<input>
<ID>IN_2</ID>169 </input>
<input>
<ID>IN_3</ID>165 </input>
<input>
<ID>IN_4</ID>173 </input>
<input>
<ID>IN_5</ID>161 </input>
<input>
<ID>IN_6</ID>167 </input>
<input>
<ID>IN_7</ID>160 </input>
<input>
<ID>IN_8</ID>170 </input>
<input>
<ID>IN_9</ID>166 </input>
<output>
<ID>OUT_0</ID>465 </output>
<output>
<ID>OUT_1</ID>467 </output>
<output>
<ID>OUT_10</ID>469 </output>
<output>
<ID>OUT_11</ID>474 </output>
<output>
<ID>OUT_12</ID>478 </output>
<output>
<ID>OUT_13</ID>470 </output>
<output>
<ID>OUT_14</ID>472 </output>
<output>
<ID>OUT_15</ID>476 </output>
<output>
<ID>OUT_2</ID>463 </output>
<output>
<ID>OUT_3</ID>464 </output>
<output>
<ID>OUT_4</ID>466 </output>
<output>
<ID>OUT_5</ID>475 </output>
<output>
<ID>OUT_6</ID>477 </output>
<output>
<ID>OUT_7</ID>468 </output>
<output>
<ID>OUT_8</ID>471 </output>
<output>
<ID>OUT_9</ID>473 </output>
<input>
<ID>clear</ID>589 </input>
<input>
<ID>clock</ID>494 </input>
<input>
<ID>count_enable</ID>587 </input>
<input>
<ID>load</ID>588 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>-10,-83</position>
<input>
<ID>IN_0</ID>497 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>36,-115</position>
<gparam>LABEL_TEXT Temporary Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>36,-63</position>
<input>
<ID>IN_0</ID>498 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>4,-136.5</position>
<gparam>LABEL_TEXT Output Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>-5,-42</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>24</ID>
<type>BX_16X1_BUS_END</type>
<position>34.5,-29.5</position>
<input>
<ID>Bus_in_0</ID>294 </input>
<input>
<ID>IN_1</ID>293 </input>
<input>
<ID>IN_10</ID>282 </input>
<input>
<ID>IN_11</ID>281 </input>
<input>
<ID>IN_2</ID>292 </input>
<input>
<ID>IN_3</ID>291 </input>
<input>
<ID>IN_4</ID>290 </input>
<input>
<ID>IN_5</ID>289 </input>
<input>
<ID>IN_6</ID>288 </input>
<input>
<ID>IN_7</ID>287 </input>
<input>
<ID>IN_8</ID>279 </input>
<input>
<ID>IN_9</ID>280 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>25</ID>
<type>BX_16X1_BUS_END</type>
<position>23,-1</position>
<input>
<ID>Bus_in_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_10</ID>13 </input>
<input>
<ID>IN_11</ID>15 </input>
<input>
<ID>IN_12</ID>10 </input>
<input>
<ID>IN_13</ID>9 </input>
<input>
<ID>IN_14</ID>12 </input>
<input>
<ID>IN_15</ID>17 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>3 </input>
<input>
<ID>IN_4</ID>4 </input>
<input>
<ID>IN_5</ID>8 </input>
<input>
<ID>IN_6</ID>5 </input>
<input>
<ID>IN_7</ID>11 </input>
<input>
<ID>IN_8</ID>16 </input>
<input>
<ID>IN_9</ID>14 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>32</ID>
<type>BB_CLOCK</type>
<position>-19,4.5</position>
<output>
<ID>CLK</ID>492 </output>
<gparam>angle 0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>33</ID>
<type>BX_16X1_BUS_END</type>
<position>24.5,-51</position>
<input>
<ID>Bus_in_0</ID>108 </input>
<input>
<ID>IN_1</ID>107 </input>
<input>
<ID>IN_10</ID>106 </input>
<input>
<ID>IN_11</ID>101 </input>
<input>
<ID>IN_2</ID>109 </input>
<input>
<ID>IN_3</ID>110 </input>
<input>
<ID>IN_4</ID>99 </input>
<input>
<ID>IN_5</ID>104 </input>
<input>
<ID>IN_6</ID>105 </input>
<input>
<ID>IN_7</ID>100 </input>
<input>
<ID>IN_8</ID>103 </input>
<input>
<ID>IN_9</ID>102 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>34</ID>
<type>BX_16X1_BUS_END</type>
<position>-13.5,-70.5</position>
<input>
<ID>Bus_in_0</ID>125 </input>
<input>
<ID>IN_1</ID>116 </input>
<input>
<ID>IN_10</ID>115 </input>
<input>
<ID>IN_11</ID>120 </input>
<input>
<ID>IN_12</ID>122 </input>
<input>
<ID>IN_13</ID>117 </input>
<input>
<ID>IN_14</ID>118 </input>
<input>
<ID>IN_15</ID>121 </input>
<input>
<ID>IN_2</ID>123 </input>
<input>
<ID>IN_3</ID>112 </input>
<input>
<ID>IN_4</ID>126 </input>
<input>
<ID>IN_5</ID>119 </input>
<input>
<ID>IN_6</ID>114 </input>
<input>
<ID>IN_7</ID>113 </input>
<input>
<ID>IN_8</ID>111 </input>
<input>
<ID>IN_9</ID>124 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>99</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>48,-55</position>
<input>
<ID>ENABLE_0</ID>693 </input>
<input>
<ID>IN_0</ID>552 </input>
<input>
<ID>IN_1</ID>557 </input>
<input>
<ID>IN_2</ID>551 </input>
<input>
<ID>IN_3</ID>556 </input>
<input>
<ID>IN_4</ID>553 </input>
<input>
<ID>IN_5</ID>554 </input>
<input>
<ID>IN_6</ID>555 </input>
<input>
<ID>IN_7</ID>558 </input>
<output>
<ID>OUT_0</ID>661 </output>
<output>
<ID>OUT_1</ID>662 </output>
<output>
<ID>OUT_2</ID>663 </output>
<output>
<ID>OUT_3</ID>664 </output>
<output>
<ID>OUT_4</ID>665 </output>
<output>
<ID>OUT_5</ID>666 </output>
<output>
<ID>OUT_6</ID>667 </output>
<output>
<ID>OUT_7</ID>668 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>100</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>52.5,-49</position>
<input>
<ID>ENABLE_0</ID>693 </input>
<input>
<ID>IN_0</ID>559 </input>
<input>
<ID>IN_1</ID>560 </input>
<input>
<ID>IN_2</ID>561 </input>
<input>
<ID>IN_3</ID>562 </input>
<output>
<ID>OUT_0</ID>657 </output>
<output>
<ID>OUT_1</ID>658 </output>
<output>
<ID>OUT_2</ID>660 </output>
<output>
<ID>OUT_3</ID>659 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>36</ID>
<type>BX_16X1_BUS_END</type>
<position>-14,-111.5</position>
<input>
<ID>Bus_in_0</ID>146 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_10</ID>147 </input>
<input>
<ID>IN_11</ID>145 </input>
<input>
<ID>IN_12</ID>152 </input>
<input>
<ID>IN_13</ID>153 </input>
<input>
<ID>IN_14</ID>155 </input>
<input>
<ID>IN_15</ID>158 </input>
<input>
<ID>IN_2</ID>150 </input>
<input>
<ID>IN_3</ID>149 </input>
<input>
<ID>IN_4</ID>148 </input>
<input>
<ID>IN_5</ID>156 </input>
<input>
<ID>IN_6</ID>143 </input>
<input>
<ID>IN_7</ID>154 </input>
<input>
<ID>IN_8</ID>151 </input>
<input>
<ID>IN_9</ID>157 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>37</ID>
<type>BX_16X1_BUS_END</type>
<position>28,-131.5</position>
<input>
<ID>Bus_in_0</ID>164 </input>
<input>
<ID>IN_1</ID>168 </input>
<input>
<ID>IN_10</ID>171 </input>
<input>
<ID>IN_11</ID>172 </input>
<input>
<ID>IN_12</ID>174 </input>
<input>
<ID>IN_13</ID>159 </input>
<input>
<ID>IN_14</ID>162 </input>
<input>
<ID>IN_15</ID>163 </input>
<input>
<ID>IN_2</ID>169 </input>
<input>
<ID>IN_3</ID>165 </input>
<input>
<ID>IN_4</ID>173 </input>
<input>
<ID>IN_5</ID>161 </input>
<input>
<ID>IN_6</ID>167 </input>
<input>
<ID>IN_7</ID>160 </input>
<input>
<ID>IN_8</ID>170 </input>
<input>
<ID>IN_9</ID>166 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>53</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>1.5,-70.5</position>
<input>
<ID>ENABLE_0</ID>694 </input>
<input>
<ID>IN_0</ID>369 </input>
<input>
<ID>IN_1</ID>374 </input>
<input>
<ID>IN_10</ID>377 </input>
<input>
<ID>IN_11</ID>379 </input>
<input>
<ID>IN_12</ID>380 </input>
<input>
<ID>IN_13</ID>381 </input>
<input>
<ID>IN_14</ID>371 </input>
<input>
<ID>IN_15</ID>382 </input>
<input>
<ID>IN_2</ID>375 </input>
<input>
<ID>IN_3</ID>367 </input>
<input>
<ID>IN_4</ID>373 </input>
<input>
<ID>IN_5</ID>372 </input>
<input>
<ID>IN_6</ID>368 </input>
<input>
<ID>IN_7</ID>378 </input>
<input>
<ID>IN_8</ID>370 </input>
<input>
<ID>IN_9</ID>376 </input>
<output>
<ID>OUT_0</ID>365 </output>
<output>
<ID>OUT_1</ID>366 </output>
<output>
<ID>OUT_10</ID>352 </output>
<output>
<ID>OUT_11</ID>357 </output>
<output>
<ID>OUT_12</ID>351 </output>
<output>
<ID>OUT_13</ID>358 </output>
<output>
<ID>OUT_14</ID>356 </output>
<output>
<ID>OUT_15</ID>359 </output>
<output>
<ID>OUT_2</ID>362 </output>
<output>
<ID>OUT_3</ID>363 </output>
<output>
<ID>OUT_4</ID>360 </output>
<output>
<ID>OUT_5</ID>361 </output>
<output>
<ID>OUT_6</ID>364 </output>
<output>
<ID>OUT_7</ID>353 </output>
<output>
<ID>OUT_8</ID>354 </output>
<output>
<ID>OUT_9</ID>355 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>54</ID>
<type>BX_16X1_BUS_END</type>
<position>6,-70.5</position>
<input>
<ID>Bus_in_0</ID>365 </input>
<input>
<ID>IN_1</ID>366 </input>
<input>
<ID>IN_10</ID>352 </input>
<input>
<ID>IN_11</ID>357 </input>
<input>
<ID>IN_12</ID>351 </input>
<input>
<ID>IN_13</ID>358 </input>
<input>
<ID>IN_14</ID>356 </input>
<input>
<ID>IN_15</ID>359 </input>
<input>
<ID>IN_2</ID>362 </input>
<input>
<ID>IN_3</ID>363 </input>
<input>
<ID>IN_4</ID>360 </input>
<input>
<ID>IN_5</ID>361 </input>
<input>
<ID>IN_6</ID>364 </input>
<input>
<ID>IN_7</ID>353 </input>
<input>
<ID>IN_8</ID>354 </input>
<input>
<ID>IN_9</ID>355 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>55</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>43.5,-90</position>
<input>
<ID>ENABLE_0</ID>695 </input>
<input>
<ID>IN_0</ID>414 </input>
<input>
<ID>IN_1</ID>399 </input>
<input>
<ID>IN_10</ID>405 </input>
<input>
<ID>IN_11</ID>403 </input>
<input>
<ID>IN_12</ID>404 </input>
<input>
<ID>IN_13</ID>406 </input>
<input>
<ID>IN_14</ID>407 </input>
<input>
<ID>IN_15</ID>409 </input>
<input>
<ID>IN_2</ID>410 </input>
<input>
<ID>IN_3</ID>400 </input>
<input>
<ID>IN_4</ID>401 </input>
<input>
<ID>IN_5</ID>408 </input>
<input>
<ID>IN_6</ID>411 </input>
<input>
<ID>IN_7</ID>412 </input>
<input>
<ID>IN_8</ID>402 </input>
<input>
<ID>IN_9</ID>413 </input>
<output>
<ID>OUT_0</ID>397 </output>
<output>
<ID>OUT_1</ID>398 </output>
<output>
<ID>OUT_10</ID>384 </output>
<output>
<ID>OUT_11</ID>389 </output>
<output>
<ID>OUT_12</ID>383 </output>
<output>
<ID>OUT_13</ID>390 </output>
<output>
<ID>OUT_14</ID>388 </output>
<output>
<ID>OUT_15</ID>391 </output>
<output>
<ID>OUT_2</ID>394 </output>
<output>
<ID>OUT_3</ID>395 </output>
<output>
<ID>OUT_4</ID>392 </output>
<output>
<ID>OUT_5</ID>393 </output>
<output>
<ID>OUT_6</ID>396 </output>
<output>
<ID>OUT_7</ID>385 </output>
<output>
<ID>OUT_8</ID>386 </output>
<output>
<ID>OUT_9</ID>387 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>56</ID>
<type>BX_16X1_BUS_END</type>
<position>48,-90</position>
<input>
<ID>Bus_in_0</ID>397 </input>
<input>
<ID>IN_1</ID>398 </input>
<input>
<ID>IN_10</ID>384 </input>
<input>
<ID>IN_11</ID>389 </input>
<input>
<ID>IN_12</ID>383 </input>
<input>
<ID>IN_13</ID>390 </input>
<input>
<ID>IN_14</ID>388 </input>
<input>
<ID>IN_15</ID>391 </input>
<input>
<ID>IN_2</ID>394 </input>
<input>
<ID>IN_3</ID>395 </input>
<input>
<ID>IN_4</ID>392 </input>
<input>
<ID>IN_5</ID>393 </input>
<input>
<ID>IN_6</ID>396 </input>
<input>
<ID>IN_7</ID>385 </input>
<input>
<ID>IN_8</ID>386 </input>
<input>
<ID>IN_9</ID>387 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>57</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>1,-111.5</position>
<input>
<ID>ENABLE_0</ID>696 </input>
<input>
<ID>IN_0</ID>431 </input>
<input>
<ID>IN_1</ID>432 </input>
<input>
<ID>IN_10</ID>439 </input>
<input>
<ID>IN_11</ID>444 </input>
<input>
<ID>IN_12</ID>443 </input>
<input>
<ID>IN_13</ID>445 </input>
<input>
<ID>IN_14</ID>442 </input>
<input>
<ID>IN_15</ID>446 </input>
<input>
<ID>IN_2</ID>433 </input>
<input>
<ID>IN_3</ID>434 </input>
<input>
<ID>IN_4</ID>435 </input>
<input>
<ID>IN_5</ID>440 </input>
<input>
<ID>IN_6</ID>441 </input>
<input>
<ID>IN_7</ID>436 </input>
<input>
<ID>IN_8</ID>437 </input>
<input>
<ID>IN_9</ID>438 </input>
<output>
<ID>OUT_0</ID>429 </output>
<output>
<ID>OUT_1</ID>430 </output>
<output>
<ID>OUT_10</ID>416 </output>
<output>
<ID>OUT_11</ID>421 </output>
<output>
<ID>OUT_12</ID>415 </output>
<output>
<ID>OUT_13</ID>422 </output>
<output>
<ID>OUT_14</ID>420 </output>
<output>
<ID>OUT_15</ID>423 </output>
<output>
<ID>OUT_2</ID>426 </output>
<output>
<ID>OUT_3</ID>427 </output>
<output>
<ID>OUT_4</ID>424 </output>
<output>
<ID>OUT_5</ID>425 </output>
<output>
<ID>OUT_6</ID>428 </output>
<output>
<ID>OUT_8</ID>418 </output>
<output>
<ID>OUT_9</ID>419 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>58</ID>
<type>BX_16X1_BUS_END</type>
<position>5.5,-111.5</position>
<input>
<ID>Bus_in_0</ID>429 </input>
<input>
<ID>IN_1</ID>430 </input>
<input>
<ID>IN_10</ID>416 </input>
<input>
<ID>IN_11</ID>421 </input>
<input>
<ID>IN_12</ID>415 </input>
<input>
<ID>IN_13</ID>422 </input>
<input>
<ID>IN_14</ID>420 </input>
<input>
<ID>IN_15</ID>423 </input>
<input>
<ID>IN_2</ID>426 </input>
<input>
<ID>IN_3</ID>427 </input>
<input>
<ID>IN_4</ID>424 </input>
<input>
<ID>IN_5</ID>425 </input>
<input>
<ID>IN_6</ID>428 </input>
<input>
<ID>IN_7</ID>417 </input>
<input>
<ID>IN_8</ID>418 </input>
<input>
<ID>IN_9</ID>419 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>59</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>43,-131.5</position>
<input>
<ID>ENABLE_0</ID>697 </input>
<input>
<ID>IN_0</ID>465 </input>
<input>
<ID>IN_1</ID>467 </input>
<input>
<ID>IN_10</ID>469 </input>
<input>
<ID>IN_11</ID>474 </input>
<input>
<ID>IN_12</ID>478 </input>
<input>
<ID>IN_13</ID>470 </input>
<input>
<ID>IN_14</ID>472 </input>
<input>
<ID>IN_15</ID>476 </input>
<input>
<ID>IN_2</ID>463 </input>
<input>
<ID>IN_3</ID>464 </input>
<input>
<ID>IN_4</ID>466 </input>
<input>
<ID>IN_5</ID>475 </input>
<input>
<ID>IN_6</ID>477 </input>
<input>
<ID>IN_7</ID>468 </input>
<input>
<ID>IN_8</ID>471 </input>
<input>
<ID>IN_9</ID>473 </input>
<output>
<ID>OUT_0</ID>461 </output>
<output>
<ID>OUT_1</ID>462 </output>
<output>
<ID>OUT_10</ID>448 </output>
<output>
<ID>OUT_11</ID>453 </output>
<output>
<ID>OUT_12</ID>447 </output>
<output>
<ID>OUT_13</ID>454 </output>
<output>
<ID>OUT_14</ID>452 </output>
<output>
<ID>OUT_15</ID>455 </output>
<output>
<ID>OUT_2</ID>458 </output>
<output>
<ID>OUT_3</ID>459 </output>
<output>
<ID>OUT_4</ID>456 </output>
<output>
<ID>OUT_5</ID>457 </output>
<output>
<ID>OUT_6</ID>460 </output>
<output>
<ID>OUT_7</ID>449 </output>
<output>
<ID>OUT_8</ID>450 </output>
<output>
<ID>OUT_9</ID>451 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>60</ID>
<type>BX_16X1_BUS_END</type>
<position>47.5,-131.5</position>
<input>
<ID>Bus_in_0</ID>461 </input>
<input>
<ID>IN_1</ID>462 </input>
<input>
<ID>IN_10</ID>448 </input>
<input>
<ID>IN_11</ID>453 </input>
<input>
<ID>IN_12</ID>447 </input>
<input>
<ID>IN_13</ID>454 </input>
<input>
<ID>IN_14</ID>452 </input>
<input>
<ID>IN_15</ID>455 </input>
<input>
<ID>IN_2</ID>458 </input>
<input>
<ID>IN_3</ID>459 </input>
<input>
<ID>IN_4</ID>456 </input>
<input>
<ID>IN_5</ID>457 </input>
<input>
<ID>IN_6</ID>460 </input>
<input>
<ID>IN_7</ID>449 </input>
<input>
<ID>IN_8</ID>450 </input>
<input>
<ID>IN_9</ID>451 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>105</ID>
<type>DA_FROM</type>
<position>44.5,13</position>
<input>
<ID>IN_0</ID>563 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID mem_w</lparam></gate>
<gate>
<ID>106</ID>
<type>DA_FROM</type>
<position>34.5,12</position>
<input>
<ID>IN_0</ID>564 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID mem_r</lparam></gate>
<gate>
<ID>107</ID>
<type>DA_FROM</type>
<position>3,-42</position>
<input>
<ID>IN_0</ID>565 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clr_addr</lparam></gate>
<gate>
<ID>108</ID>
<type>DA_FROM</type>
<position>-4.5,-22.5</position>
<input>
<ID>IN_0</ID>566 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_addr</lparam></gate>
<gate>
<ID>111</ID>
<type>DA_FROM</type>
<position>2,-20.5</position>
<input>
<ID>IN_0</ID>568 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID inc_addr</lparam></gate>
<gate>
<ID>112</ID>
<type>DA_FROM</type>
<position>44,-63</position>
<input>
<ID>IN_0</ID>569 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clr_pc</lparam></gate>
<gate>
<ID>113</ID>
<type>DA_FROM</type>
<position>35,-44</position>
<input>
<ID>IN_0</ID>570 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_pc</lparam></gate>
<gate>
<ID>114</ID>
<type>DA_FROM</type>
<position>44,-43</position>
<input>
<ID>IN_0</ID>572 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID inc_pc</lparam></gate>
<gate>
<ID>115</ID>
<type>EE_VDD</type>
<position>41,-44</position>
<output>
<ID>OUT_0</ID>571 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>116</ID>
<type>DA_FROM</type>
<position>-2,-83</position>
<input>
<ID>IN_0</ID>573 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clr_data</lparam></gate>
<gate>
<ID>117</ID>
<type>DA_FROM</type>
<position>-3,-57.5</position>
<input>
<ID>IN_0</ID>575 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID inc_dr</lparam></gate>
<gate>
<ID>118</ID>
<type>EE_VDD</type>
<position>-5,-59.5</position>
<output>
<ID>OUT_0</ID>574 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>119</ID>
<type>DA_FROM</type>
<position>-10.5,-59.5</position>
<input>
<ID>IN_0</ID>576 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_dr</lparam></gate>
<gate>
<ID>120</ID>
<type>DA_FROM</type>
<position>38.5,-77</position>
<input>
<ID>IN_0</ID>577 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID inc_ac</lparam></gate>
<gate>
<ID>121</ID>
<type>EE_VDD</type>
<position>37,-79</position>
<output>
<ID>OUT_0</ID>578 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>122</ID>
<type>EE_VDD</type>
<position>-5.5,-100.5</position>
<output>
<ID>OUT_0</ID>579 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>124</ID>
<type>EE_VDD</type>
<position>4.5,-141</position>
<output>
<ID>OUT_0</ID>581 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>31,-79</position>
<input>
<ID>IN_0</ID>582 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_ac</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>40,-102.5</position>
<input>
<ID>IN_0</ID>583 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clr_ac</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>-10.5,-101</position>
<input>
<ID>IN_0</ID>585 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_ir</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>38.5,-118</position>
<input>
<ID>IN_0</ID>587 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID inc_tr</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>31,-120.5</position>
<input>
<ID>IN_0</ID>588 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_tr</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>39.5,-144.5</position>
<input>
<ID>IN_0</ID>589 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clr_tr</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>0,-141</position>
<input>
<ID>IN_0</ID>591 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ld_or</lparam></gate>
<gate>
<ID>136</ID>
<type>BX_16X1_BUS_END</type>
<position>-11.5,-144</position>
<input>
<ID>Bus_in_0</ID>609 </input>
<input>
<ID>IN_1</ID>610 </input>
<input>
<ID>IN_2</ID>611 </input>
<input>
<ID>IN_3</ID>614 </input>
<input>
<ID>IN_4</ID>615 </input>
<input>
<ID>IN_5</ID>616 </input>
<input>
<ID>IN_6</ID>612 </input>
<input>
<ID>IN_7</ID>613 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>137</ID>
<type>BX_16X1_BUS_END</type>
<position>61.5,-51</position>
<input>
<ID>Bus_in_0</ID>661 </input>
<input>
<ID>IN_1</ID>662 </input>
<input>
<ID>IN_10</ID>660 </input>
<input>
<ID>IN_11</ID>659 </input>
<input>
<ID>IN_2</ID>663 </input>
<input>
<ID>IN_3</ID>664 </input>
<input>
<ID>IN_4</ID>665 </input>
<input>
<ID>IN_5</ID>666 </input>
<input>
<ID>IN_6</ID>667 </input>
<input>
<ID>IN_7</ID>668 </input>
<input>
<ID>IN_8</ID>657 </input>
<input>
<ID>IN_9</ID>658 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>164</ID>
<type>DA_FROM</type>
<position>55.5,-40</position>
<input>
<ID>IN_0</ID>693 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_pc</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>8,-59.5</position>
<input>
<ID>IN_0</ID>694 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_dr</lparam></gate>
<gate>
<ID>166</ID>
<type>DA_FROM</type>
<position>51.5,-79</position>
<input>
<ID>IN_0</ID>695 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_ac</lparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>7,-100.5</position>
<input>
<ID>IN_0</ID>696 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_ir</lparam></gate>
<gate>
<ID>168</ID>
<type>DA_FROM</type>
<position>48,-119.5</position>
<input>
<ID>IN_0</ID>697 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_tr</lparam></gate>
<gate>
<ID>27</ID>
<type>BX_16X1_BUS_END</type>
<position>-15.5,-29.5</position>
<input>
<ID>Bus_in_0</ID>95 </input>
<input>
<ID>IN_1</ID>179 </input>
<input>
<ID>IN_10</ID>177 </input>
<input>
<ID>IN_11</ID>178 </input>
<input>
<ID>IN_2</ID>93 </input>
<input>
<ID>IN_3</ID>96 </input>
<input>
<ID>IN_4</ID>97 </input>
<input>
<ID>IN_5</ID>98 </input>
<input>
<ID>IN_6</ID>176 </input>
<input>
<ID>IN_7</ID>94 </input>
<input>
<ID>IN_8</ID>180 </input>
<input>
<ID>IN_9</ID>175 </input>
<input>
<ID>OUT</ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>66</ID>
<type>BX_16X1_BUS_END</type>
<position>9,-29.5</position>
<input>
<ID>Bus_in_0</ID>188 </input>
<input>
<ID>IN_1</ID>182 </input>
<input>
<ID>IN_10</ID>191 </input>
<input>
<ID>IN_11</ID>192 </input>
<input>
<ID>IN_2</ID>190 </input>
<input>
<ID>IN_3</ID>189 </input>
<input>
<ID>IN_4</ID>181 </input>
<input>
<ID>IN_5</ID>183 </input>
<input>
<ID>IN_6</ID>184 </input>
<input>
<ID>IN_7</ID>185 </input>
<input>
<ID>IN_8</ID>187 </input>
<input>
<ID>IN_9</ID>186 </input>
<input>
<ID>OUT</ID>205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>67</ID>
<type>BX_16X1_BUS_END</type>
<position>10.5,14.5</position>
<input>
<ID>Bus_in_0</ID>197 </input>
<input>
<ID>IN_1</ID>198 </input>
<input>
<ID>IN_10</ID>203 </input>
<input>
<ID>IN_11</ID>204 </input>
<input>
<ID>IN_2</ID>195 </input>
<input>
<ID>IN_3</ID>201 </input>
<input>
<ID>IN_4</ID>199 </input>
<input>
<ID>IN_5</ID>202 </input>
<input>
<ID>IN_6</ID>200 </input>
<input>
<ID>IN_7</ID>193 </input>
<input>
<ID>IN_8</ID>194 </input>
<input>
<ID>IN_9</ID>196 </input>
<input>
<ID>OUT</ID>205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>68</ID>
<type>BX_16X1_BUS_END</type>
<position>20.5,-29.5</position>
<input>
<ID>Bus_in_0</ID>272 </input>
<input>
<ID>IN_1</ID>276 </input>
<input>
<ID>IN_10</ID>285 </input>
<input>
<ID>IN_11</ID>286 </input>
<input>
<ID>IN_2</ID>273 </input>
<input>
<ID>IN_3</ID>275 </input>
<input>
<ID>IN_4</ID>277 </input>
<input>
<ID>IN_5</ID>271 </input>
<input>
<ID>IN_6</ID>274 </input>
<input>
<ID>IN_7</ID>278 </input>
<input>
<ID>IN_8</ID>283 </input>
<input>
<ID>IN_9</ID>284 </input>
<input>
<ID>OUT</ID>205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>33,-18</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID bus_ar</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>28.5,-97.5</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc0</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>19.5,-96.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc1</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>28.5,-95.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc2</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>19.5,-94.5</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc3</lparam></gate>
<gate>
<ID>85</ID>
<type>DA_FROM</type>
<position>28.5,-93.5</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc4</lparam></gate>
<gate>
<ID>86</ID>
<type>DA_FROM</type>
<position>19.5,-92.5</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc5</lparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>28.5,-91.5</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc6</lparam></gate>
<gate>
<ID>88</ID>
<type>DA_FROM</type>
<position>19.5,-90.5</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc7</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>28.5,-89.5</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc8</lparam></gate>
<gate>
<ID>90</ID>
<type>DA_FROM</type>
<position>19.5,-88.5</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc9</lparam></gate>
<gate>
<ID>91</ID>
<type>DA_FROM</type>
<position>28.5,-87.5</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc10</lparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>19.5,-86.5</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc11</lparam></gate>
<gate>
<ID>93</ID>
<type>DA_FROM</type>
<position>28.5,-85.5</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc12</lparam></gate>
<gate>
<ID>94</ID>
<type>DA_FROM</type>
<position>19.5,-84.5</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc13</lparam></gate>
<gate>
<ID>95</ID>
<type>DA_FROM</type>
<position>28.5,-83.5</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc14</lparam></gate>
<gate>
<ID>96</ID>
<type>DA_FROM</type>
<position>19.5,-82.5</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID acc15</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>-60.5,20.5</position>
<gparam>LABEL_TEXT Mano Machine</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>-52,14</position>
<gparam>LABEL_TEXT Checkpoint 1 - Brandon Aikman</gparam>
<gparam>TEXT_HEIGHT 2.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>25.5,-33.5</position>
<input>
<ID>ENABLE_0</ID>295 </input>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>276 </input>
<input>
<ID>IN_2</ID>273 </input>
<input>
<ID>IN_3</ID>275 </input>
<input>
<ID>IN_4</ID>277 </input>
<input>
<ID>IN_5</ID>271 </input>
<input>
<ID>IN_6</ID>274 </input>
<input>
<ID>IN_7</ID>278 </input>
<output>
<ID>OUT_0</ID>294 </output>
<output>
<ID>OUT_1</ID>293 </output>
<output>
<ID>OUT_2</ID>292 </output>
<output>
<ID>OUT_3</ID>291 </output>
<output>
<ID>OUT_4</ID>290 </output>
<output>
<ID>OUT_5</ID>289 </output>
<output>
<ID>OUT_6</ID>288 </output>
<output>
<ID>OUT_7</ID>287 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>102</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>30,-27.5</position>
<input>
<ID>ENABLE_0</ID>295 </input>
<input>
<ID>IN_0</ID>283 </input>
<input>
<ID>IN_1</ID>284 </input>
<input>
<ID>IN_2</ID>285 </input>
<input>
<ID>IN_3</ID>286 </input>
<output>
<ID>OUT_0</ID>279 </output>
<output>
<ID>OUT_1</ID>280 </output>
<output>
<ID>OUT_2</ID>282 </output>
<output>
<ID>OUT_3</ID>281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>4 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,1,26.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_4</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>25</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>491 </ID>
<shape>
<hsegment>
<ID>8</ID>
<points>32,14,32.5,14</points>
<connection>
<GID>2</GID>
<name>write_clock</name></connection>
<connection>
<GID>74</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,1,16.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_14</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_14</name></connection>
<connection>
<GID>25</GID>
<name>IN_14</name></connection></vsegment></shape></wire>
<wire>
<ID>570 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-45.5,39,-44</points>
<connection>
<GID>12</GID>
<name>load</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-44,39,-44</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>112 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-75,-11,-75</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<connection>
<GID>34</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>15 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,1,19.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_11</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_11</name></connection>
<connection>
<GID>25</GID>
<name>IN_11</name></connection></vsegment></shape></wire>
<wire>
<ID>657 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-50.5,59.5,-50.5</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<connection>
<GID>137</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>560 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-49.5,50.5,-49.5</points>
<connection>
<GID>12</GID>
<name>OUT_9</name></connection>
<connection>
<GID>100</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>122 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-66,-11,-66</points>
<connection>
<GID>8</GID>
<name>IN_12</name></connection>
<connection>
<GID>34</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>2 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,1,28.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_2</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>25</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>9 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,1,17.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_13</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_13</name></connection>
<connection>
<GID>25</GID>
<name>IN_13</name></connection></vsegment></shape></wire>
<wire>
<ID>17 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,1,15.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_15</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_15</name></connection>
<connection>
<GID>25</GID>
<name>IN_15</name></connection></vsegment></shape></wire>
<wire>
<ID>3 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,1,27.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_3</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>25</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>661 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-58.5,59.5,-58.5</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<connection>
<GID>137</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>564 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,12,32.5,12</points>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>126 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-74,-11,-74</points>
<connection>
<GID>8</GID>
<name>IN_4</name></connection>
<connection>
<GID>34</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>422 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-106,3.5,-106</points>
<connection>
<GID>57</GID>
<name>OUT_13</name></connection>
<connection>
<GID>58</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>571 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-45.5,41,-45</points>
<connection>
<GID>12</GID>
<name>count_up</name></connection>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,1,20.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_10</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_10</name></connection>
<connection>
<GID>25</GID>
<name>IN_10</name></connection></vsegment></shape></wire>
<wire>
<ID>120 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-67,-11,-67</points>
<connection>
<GID>8</GID>
<name>IN_11</name></connection>
<connection>
<GID>34</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>665 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-54.5,59.5,-54.5</points>
<connection>
<GID>99</GID>
<name>OUT_4</name></connection>
<connection>
<GID>137</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>572 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-45.5,40,-43</points>
<connection>
<GID>12</GID>
<name>count_enable</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-43,42,-43</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>493 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-158,2.5,-153.5</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<intersection>-158 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-158,2.5,-158</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,1,30.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_0</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>Bus_in_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,1,29.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_1</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>25</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>497 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-83,-7,-80</points>
<connection>
<GID>8</GID>
<name>clock</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,-83,-7,-83</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>10 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,1,18.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_12</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_12</name></connection>
<connection>
<GID>25</GID>
<name>IN_12</name></connection></vsegment></shape></wire>
<wire>
<ID>8 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,1,25.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_5</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>25</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>414 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-97.5,41.5,-97.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>563 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,13,42.5,13</points>
<connection>
<GID>2</GID>
<name>write_enable</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,1,24.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_6</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>25</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>492 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-15,4.5,-9,4.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>11 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,1,23.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_7</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>25</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>16 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,1,22.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_8</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_8</name></connection>
<connection>
<GID>25</GID>
<name>IN_8</name></connection></vsegment></shape></wire>
<wire>
<ID>14 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,1,21.5,1.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_9</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_9</name></connection>
<connection>
<GID>25</GID>
<name>IN_9</name></connection></vsegment></shape></wire>
<wire>
<ID>459 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-136,45.5,-136</points>
<connection>
<GID>59</GID>
<name>OUT_3</name></connection>
<connection>
<GID>60</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>108 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-58.5,35,-58.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>33</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>107 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-57.5,35,-57.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<connection>
<GID>33</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>465 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-139,41,-139</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>106 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-48.5,35,-48.5</points>
<connection>
<GID>12</GID>
<name>IN_10</name></connection>
<connection>
<GID>33</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>101 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-47.5,35,-47.5</points>
<connection>
<GID>12</GID>
<name>IN_11</name></connection>
<connection>
<GID>33</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>109 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-56.5,35,-56.5</points>
<connection>
<GID>12</GID>
<name>IN_2</name></connection>
<connection>
<GID>33</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>469 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-129,41,-129</points>
<connection>
<GID>18</GID>
<name>OUT_10</name></connection>
<connection>
<GID>59</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>110 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-55.5,35,-55.5</points>
<connection>
<GID>12</GID>
<name>IN_3</name></connection>
<connection>
<GID>33</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>99 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-54.5,35,-54.5</points>
<connection>
<GID>12</GID>
<name>IN_4</name></connection>
<connection>
<GID>33</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>562 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-47.5,50.5,-47.5</points>
<connection>
<GID>12</GID>
<name>OUT_11</name></connection>
<connection>
<GID>100</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>471 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-131,41,-131</points>
<connection>
<GID>18</GID>
<name>OUT_8</name></connection>
<connection>
<GID>59</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>104 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-53.5,35,-53.5</points>
<connection>
<GID>12</GID>
<name>IN_5</name></connection>
<connection>
<GID>33</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>386 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-89.5,46,-89.5</points>
<connection>
<GID>55</GID>
<name>OUT_8</name></connection>
<connection>
<GID>56</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>551 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-56.5,46,-56.5</points>
<connection>
<GID>12</GID>
<name>OUT_2</name></connection>
<connection>
<GID>99</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>105 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-52.5,35,-52.5</points>
<connection>
<GID>12</GID>
<name>IN_6</name></connection>
<connection>
<GID>33</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>558 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-51.5,46,-51.5</points>
<connection>
<GID>12</GID>
<name>OUT_7</name></connection>
<connection>
<GID>99</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>451 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-130,45.5,-130</points>
<connection>
<GID>59</GID>
<name>OUT_9</name></connection>
<connection>
<GID>60</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>100 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-51.5,35,-51.5</points>
<connection>
<GID>12</GID>
<name>IN_7</name></connection>
<connection>
<GID>33</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>376 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-69,-0.5,-69</points>
<connection>
<GID>8</GID>
<name>OUT_9</name></connection>
<connection>
<GID>53</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>553 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-54.5,46,-54.5</points>
<connection>
<GID>12</GID>
<name>OUT_4</name></connection>
<connection>
<GID>99</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>103 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-50.5,35,-50.5</points>
<connection>
<GID>12</GID>
<name>IN_8</name></connection>
<connection>
<GID>33</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>461 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-139,45.5,-139</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<connection>
<GID>60</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>102 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-49.5,35,-49.5</points>
<connection>
<GID>12</GID>
<name>IN_9</name></connection>
<connection>
<GID>33</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>264 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-82.5,31,-82.5</points>
<connection>
<GID>14</GID>
<name>IN_15</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>569 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-63,41,-60.5</points>
<connection>
<GID>12</GID>
<name>clear</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-63,42,-63</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>498 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-63,39,-60.5</points>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-63,39,-63</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>552 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-58.5,46,-58.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>380 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-66,-0.5,-66</points>
<connection>
<GID>8</GID>
<name>OUT_12</name></connection>
<connection>
<GID>53</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>557 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-57.5,46,-57.5</points>
<connection>
<GID>12</GID>
<name>OUT_1</name></connection>
<connection>
<GID>99</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>256 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-95.5,31,-95.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<connection>
<GID>75</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>561 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-48.5,50.5,-48.5</points>
<connection>
<GID>12</GID>
<name>OUT_10</name></connection>
<connection>
<GID>100</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>556 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-55.5,46,-55.5</points>
<connection>
<GID>12</GID>
<name>OUT_3</name></connection>
<connection>
<GID>99</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>554 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-53.5,46,-53.5</points>
<connection>
<GID>12</GID>
<name>OUT_5</name></connection>
<connection>
<GID>99</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>406 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-84.5,41.5,-84.5</points>
<connection>
<GID>14</GID>
<name>OUT_13</name></connection>
<connection>
<GID>55</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>555 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-52.5,46,-52.5</points>
<connection>
<GID>12</GID>
<name>OUT_6</name></connection>
<connection>
<GID>99</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>394 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-95.5,46,-95.5</points>
<connection>
<GID>55</GID>
<name>OUT_2</name></connection>
<connection>
<GID>56</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>559 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-50.5,50.5,-50.5</points>
<connection>
<GID>12</GID>
<name>OUT_8</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>432 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-118,-1,-118</points>
<connection>
<GID>16</GID>
<name>OUT_1</name></connection>
<connection>
<GID>57</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>609 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-151.5,-0.5,-151.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>136</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>610 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-150.5,-0.5,-150.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>136</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>462 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-138,45.5,-138</points>
<connection>
<GID>59</GID>
<name>OUT_1</name></connection>
<connection>
<GID>60</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>611 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-149.5,-0.5,-149.5</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<connection>
<GID>136</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>614 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-148.5,-0.5,-148.5</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<connection>
<GID>136</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>450 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-131,45.5,-131</points>
<connection>
<GID>59</GID>
<name>OUT_8</name></connection>
<connection>
<GID>60</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>615 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-147.5,-0.5,-147.5</points>
<connection>
<GID>4</GID>
<name>IN_4</name></connection>
<connection>
<GID>136</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>281 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32,-26,32.5,-26</points>
<connection>
<GID>102</GID>
<name>OUT_3</name></connection>
<connection>
<GID>24</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>616 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-146.5,-0.5,-146.5</points>
<connection>
<GID>4</GID>
<name>IN_5</name></connection>
<connection>
<GID>136</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>277 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-33,23.5,-33</points>
<connection>
<GID>68</GID>
<name>IN_4</name></connection>
<connection>
<GID>101</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>612 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-145.5,-0.5,-145.5</points>
<connection>
<GID>4</GID>
<name>IN_6</name></connection>
<connection>
<GID>136</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>436 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-112,-1,-112</points>
<connection>
<GID>16</GID>
<name>OUT_7</name></connection>
<connection>
<GID>57</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>613 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-144.5,-0.5,-144.5</points>
<connection>
<GID>4</GID>
<name>IN_7</name></connection>
<connection>
<GID>136</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>404 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-85.5,41.5,-85.5</points>
<connection>
<GID>14</GID>
<name>OUT_12</name></connection>
<connection>
<GID>55</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>581 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-142.5,4.5,-142</points>
<connection>
<GID>4</GID>
<name>count_up</name></connection>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>591 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-142.5,2.5,-141</points>
<connection>
<GID>4</GID>
<name>load</name></connection>
<intersection>-141 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-141,2.5,-141</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>583 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-102.5,37,-99.5</points>
<connection>
<GID>14</GID>
<name>clear</name></connection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-102.5,38,-102.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>496 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-102.5,35,-99.5</points>
<connection>
<GID>14</GID>
<name>clock</name></connection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-102.5,35,-102.5</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>400 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-94.5,41.5,-94.5</points>
<connection>
<GID>14</GID>
<name>OUT_3</name></connection>
<connection>
<GID>55</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>577 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-80.5,36,-77</points>
<connection>
<GID>14</GID>
<name>count_enable</name></connection>
<intersection>-77 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-77,36.5,-77</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>578 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-80.5,37,-80</points>
<connection>
<GID>14</GID>
<name>count_up</name></connection>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>582 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-80.5,35,-79</points>
<connection>
<GID>14</GID>
<name>load</name></connection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-79,35,-79</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>399 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-96.5,41.5,-96.5</points>
<connection>
<GID>14</GID>
<name>OUT_1</name></connection>
<connection>
<GID>55</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>405 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-87.5,41.5,-87.5</points>
<connection>
<GID>14</GID>
<name>OUT_10</name></connection>
<connection>
<GID>55</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>403 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-86.5,41.5,-86.5</points>
<connection>
<GID>14</GID>
<name>OUT_11</name></connection>
<connection>
<GID>55</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>407 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-83.5,41.5,-83.5</points>
<connection>
<GID>14</GID>
<name>OUT_14</name></connection>
<connection>
<GID>55</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>409 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-82.5,41.5,-82.5</points>
<connection>
<GID>14</GID>
<name>OUT_15</name></connection>
<connection>
<GID>55</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>575 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-61,-6,-57.5</points>
<connection>
<GID>8</GID>
<name>count_enable</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-57.5,-5,-57.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>410 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-95.5,41.5,-95.5</points>
<connection>
<GID>14</GID>
<name>OUT_2</name></connection>
<connection>
<GID>55</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>401 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-93.5,41.5,-93.5</points>
<connection>
<GID>14</GID>
<name>OUT_4</name></connection>
<connection>
<GID>55</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>585 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-102,-7.5,-101</points>
<connection>
<GID>16</GID>
<name>load</name></connection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-101,-7.5,-101</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>408 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-92.5,41.5,-92.5</points>
<connection>
<GID>14</GID>
<name>OUT_5</name></connection>
<connection>
<GID>55</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>411 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-91.5,41.5,-91.5</points>
<connection>
<GID>14</GID>
<name>OUT_6</name></connection>
<connection>
<GID>55</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>589 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-144.5,36.5,-141</points>
<connection>
<GID>18</GID>
<name>clear</name></connection>
<intersection>-144.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-144.5,37.5,-144.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>412 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-90.5,41.5,-90.5</points>
<connection>
<GID>14</GID>
<name>OUT_7</name></connection>
<connection>
<GID>55</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>402 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-89.5,41.5,-89.5</points>
<connection>
<GID>14</GID>
<name>OUT_8</name></connection>
<connection>
<GID>55</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>413 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-88.5,41.5,-88.5</points>
<connection>
<GID>14</GID>
<name>OUT_9</name></connection>
<connection>
<GID>55</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>415 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-107,3.5,-107</points>
<connection>
<GID>57</GID>
<name>OUT_12</name></connection>
<connection>
<GID>58</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>423 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-104,3.5,-104</points>
<connection>
<GID>57</GID>
<name>OUT_15</name></connection>
<connection>
<GID>58</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>260 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-89.5,31,-89.5</points>
<connection>
<GID>14</GID>
<name>IN_8</name></connection>
<connection>
<GID>89</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>565 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-42,0,-39</points>
<connection>
<GID>6</GID>
<name>clear</name></connection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>0,-42,1,-42</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>499 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-42,-2,-39</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3,-42,-2,-42</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>568 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-24,-1,-20.5</points>
<connection>
<GID>6</GID>
<name>count_enable</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1,-20.5,0,-20.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>566 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-24,-2,-22.5</points>
<connection>
<GID>6</GID>
<name>load</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-22.5,-2,-22.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>352 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-68,4,-68</points>
<connection>
<GID>53</GID>
<name>OUT_10</name></connection>
<connection>
<GID>54</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>360 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-74,4,-74</points>
<connection>
<GID>53</GID>
<name>OUT_4</name></connection>
<connection>
<GID>54</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>195 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,9,14,9</points>
<connection>
<GID>2</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>67</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>356 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-64,4,-64</points>
<connection>
<GID>53</GID>
<name>OUT_14</name></connection>
<connection>
<GID>54</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>125 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-78,-11,-78</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>467 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-138,41,-138</points>
<connection>
<GID>18</GID>
<name>OUT_1</name></connection>
<connection>
<GID>59</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>116 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-77,-11,-77</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>115 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-68,-11,-68</points>
<connection>
<GID>8</GID>
<name>IN_10</name></connection>
<connection>
<GID>34</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>117 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-65,-11,-65</points>
<connection>
<GID>8</GID>
<name>IN_13</name></connection>
<connection>
<GID>34</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>477 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-133,41,-133</points>
<connection>
<GID>18</GID>
<name>OUT_6</name></connection>
<connection>
<GID>59</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>118 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-64,-11,-64</points>
<connection>
<GID>8</GID>
<name>IN_14</name></connection>
<connection>
<GID>34</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>121 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-63,-11,-63</points>
<connection>
<GID>8</GID>
<name>IN_15</name></connection>
<connection>
<GID>34</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>123 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-76,-11,-76</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<connection>
<GID>34</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>119 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-73,-11,-73</points>
<connection>
<GID>8</GID>
<name>IN_5</name></connection>
<connection>
<GID>34</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>473 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-130,41,-130</points>
<connection>
<GID>18</GID>
<name>OUT_9</name></connection>
<connection>
<GID>59</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>114 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-72,-11,-72</points>
<connection>
<GID>8</GID>
<name>IN_6</name></connection>
<connection>
<GID>34</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>113 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-71,-11,-71</points>
<connection>
<GID>8</GID>
<name>IN_7</name></connection>
<connection>
<GID>34</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>111 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-70,-11,-70</points>
<connection>
<GID>8</GID>
<name>IN_8</name></connection>
<connection>
<GID>34</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>475 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-134,41,-134</points>
<connection>
<GID>18</GID>
<name>OUT_5</name></connection>
<connection>
<GID>59</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>124 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-69,-11,-69</points>
<connection>
<GID>8</GID>
<name>IN_9</name></connection>
<connection>
<GID>34</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>268 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-90.5,31,-90.5</points>
<connection>
<GID>14</GID>
<name>IN_7</name></connection>
<connection>
<GID>88</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>573 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-83,-5,-80</points>
<connection>
<GID>8</GID>
<name>clear</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-83,-4,-83</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>574 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-61,-5,-60.5</points>
<connection>
<GID>8</GID>
<name>count_up</name></connection>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>369 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-78,-0.5,-78</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>53</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>576 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-61,-7,-59.5</points>
<connection>
<GID>8</GID>
<name>load</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-59.5,-7,-59.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>374 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-77,-0.5,-77</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<connection>
<GID>53</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>377 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-68,-0.5,-68</points>
<connection>
<GID>8</GID>
<name>OUT_10</name></connection>
<connection>
<GID>53</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>379 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-67,-0.5,-67</points>
<connection>
<GID>8</GID>
<name>OUT_11</name></connection>
<connection>
<GID>53</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>588 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-122,34.5,-120.5</points>
<connection>
<GID>18</GID>
<name>load</name></connection>
<intersection>-120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-120.5,34.5,-120.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>381 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-65,-0.5,-65</points>
<connection>
<GID>8</GID>
<name>OUT_13</name></connection>
<connection>
<GID>53</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>371 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-64,-0.5,-64</points>
<connection>
<GID>8</GID>
<name>OUT_14</name></connection>
<connection>
<GID>53</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>382 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-63,-0.5,-63</points>
<connection>
<GID>8</GID>
<name>OUT_15</name></connection>
<connection>
<GID>53</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>375 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-76,-0.5,-76</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<connection>
<GID>53</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>367 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-75,-0.5,-75</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<connection>
<GID>53</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>373 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-74,-0.5,-74</points>
<connection>
<GID>8</GID>
<name>OUT_4</name></connection>
<connection>
<GID>53</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>372 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-73,-0.5,-73</points>
<connection>
<GID>8</GID>
<name>OUT_5</name></connection>
<connection>
<GID>53</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>368 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-72,-0.5,-72</points>
<connection>
<GID>8</GID>
<name>OUT_6</name></connection>
<connection>
<GID>53</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>378 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-71,-0.5,-71</points>
<connection>
<GID>8</GID>
<name>OUT_7</name></connection>
<connection>
<GID>53</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>370 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-70,-0.5,-70</points>
<connection>
<GID>8</GID>
<name>OUT_8</name></connection>
<connection>
<GID>53</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>494 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-144.5,34.5,-141</points>
<connection>
<GID>18</GID>
<name>clock</name></connection>
<intersection>-144.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-144.5,34.5,-144.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>495 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-124.5,-7.5,-121</points>
<connection>
<GID>16</GID>
<name>clock</name></connection>
<intersection>-124.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,-124.5,-7.5,-124.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>146 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-119,-11.5,-119</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>144 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-118,-11.5,-118</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<connection>
<GID>36</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>147 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-109,-11.5,-109</points>
<connection>
<GID>16</GID>
<name>IN_10</name></connection>
<connection>
<GID>36</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>145 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-108,-11.5,-108</points>
<connection>
<GID>16</GID>
<name>IN_11</name></connection>
<connection>
<GID>36</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>152 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-107,-11.5,-107</points>
<connection>
<GID>16</GID>
<name>IN_12</name></connection>
<connection>
<GID>36</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>153 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-106,-11.5,-106</points>
<connection>
<GID>16</GID>
<name>IN_13</name></connection>
<connection>
<GID>36</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>155 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-105,-11.5,-105</points>
<connection>
<GID>16</GID>
<name>IN_14</name></connection>
<connection>
<GID>36</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>158 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-104,-11.5,-104</points>
<connection>
<GID>16</GID>
<name>IN_15</name></connection>
<connection>
<GID>36</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>150 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-117,-11.5,-117</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<connection>
<GID>36</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>149 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-116,-11.5,-116</points>
<connection>
<GID>16</GID>
<name>IN_3</name></connection>
<connection>
<GID>36</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>148 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-115,-11.5,-115</points>
<connection>
<GID>16</GID>
<name>IN_4</name></connection>
<connection>
<GID>36</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>156 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-114,-11.5,-114</points>
<connection>
<GID>16</GID>
<name>IN_5</name></connection>
<connection>
<GID>36</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>288 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-31,32.5,-31</points>
<connection>
<GID>101</GID>
<name>OUT_6</name></connection>
<connection>
<GID>24</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>143 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-113,-11.5,-113</points>
<connection>
<GID>16</GID>
<name>IN_6</name></connection>
<connection>
<GID>36</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>154 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-112,-11.5,-112</points>
<connection>
<GID>16</GID>
<name>IN_7</name></connection>
<connection>
<GID>36</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>151 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-111,-11.5,-111</points>
<connection>
<GID>16</GID>
<name>IN_8</name></connection>
<connection>
<GID>36</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>157 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-110,-11.5,-110</points>
<connection>
<GID>16</GID>
<name>IN_9</name></connection>
<connection>
<GID>36</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>579 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>-5.5,-102,-5.5,-101.5</points>
<connection>
<GID>16</GID>
<name>count_up</name></connection>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>431 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-119,-1,-119</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>439 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-109,-1,-109</points>
<connection>
<GID>16</GID>
<name>OUT_10</name></connection>
<connection>
<GID>57</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>444 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-108,-1,-108</points>
<connection>
<GID>16</GID>
<name>OUT_11</name></connection>
<connection>
<GID>57</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>443 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-107,-1,-107</points>
<connection>
<GID>16</GID>
<name>OUT_12</name></connection>
<connection>
<GID>57</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>445 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-106,-1,-106</points>
<connection>
<GID>16</GID>
<name>OUT_13</name></connection>
<connection>
<GID>57</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>442 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-105,-1,-105</points>
<connection>
<GID>16</GID>
<name>OUT_14</name></connection>
<connection>
<GID>57</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>446 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-104,-1,-104</points>
<connection>
<GID>16</GID>
<name>OUT_15</name></connection>
<connection>
<GID>57</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>433 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-117,-1,-117</points>
<connection>
<GID>16</GID>
<name>OUT_2</name></connection>
<connection>
<GID>57</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>434 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-116,-1,-116</points>
<connection>
<GID>16</GID>
<name>OUT_3</name></connection>
<connection>
<GID>57</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>435 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-115,-1,-115</points>
<connection>
<GID>16</GID>
<name>OUT_4</name></connection>
<connection>
<GID>57</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>440 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-114,-1,-114</points>
<connection>
<GID>16</GID>
<name>OUT_5</name></connection>
<connection>
<GID>57</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>441 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-113,-1,-113</points>
<connection>
<GID>16</GID>
<name>OUT_6</name></connection>
<connection>
<GID>57</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>437 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-111,-1,-111</points>
<connection>
<GID>16</GID>
<name>OUT_8</name></connection>
<connection>
<GID>57</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>438 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-1.5,-110,-1,-110</points>
<connection>
<GID>16</GID>
<name>OUT_9</name></connection>
<connection>
<GID>57</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>164 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-139,30.5,-139</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>37</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>168 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-138,30.5,-138</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<connection>
<GID>37</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>171 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-129,30.5,-129</points>
<connection>
<GID>18</GID>
<name>IN_10</name></connection>
<connection>
<GID>37</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>172 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-128,30.5,-128</points>
<connection>
<GID>18</GID>
<name>IN_11</name></connection>
<connection>
<GID>37</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>174 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-127,30.5,-127</points>
<connection>
<GID>18</GID>
<name>IN_12</name></connection>
<connection>
<GID>37</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>159 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-126,30.5,-126</points>
<connection>
<GID>18</GID>
<name>IN_13</name></connection>
<connection>
<GID>37</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>162 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-125,30.5,-125</points>
<connection>
<GID>18</GID>
<name>IN_14</name></connection>
<connection>
<GID>37</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>163 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-124,30.5,-124</points>
<connection>
<GID>18</GID>
<name>IN_15</name></connection>
<connection>
<GID>37</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>169 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-137,30.5,-137</points>
<connection>
<GID>18</GID>
<name>IN_2</name></connection>
<connection>
<GID>37</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>165 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-136,30.5,-136</points>
<connection>
<GID>18</GID>
<name>IN_3</name></connection>
<connection>
<GID>37</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>173 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-135,30.5,-135</points>
<connection>
<GID>18</GID>
<name>IN_4</name></connection>
<connection>
<GID>37</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>161 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-134,30.5,-134</points>
<connection>
<GID>18</GID>
<name>IN_5</name></connection>
<connection>
<GID>37</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>167 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-133,30.5,-133</points>
<connection>
<GID>18</GID>
<name>IN_6</name></connection>
<connection>
<GID>37</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>160 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-132,30.5,-132</points>
<connection>
<GID>18</GID>
<name>IN_7</name></connection>
<connection>
<GID>37</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>170 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-131,30.5,-131</points>
<connection>
<GID>18</GID>
<name>IN_8</name></connection>
<connection>
<GID>37</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>166 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30,-130,30.5,-130</points>
<connection>
<GID>18</GID>
<name>IN_9</name></connection>
<connection>
<GID>37</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>587 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-122,35.5,-118</points>
<connection>
<GID>18</GID>
<name>count_enable</name></connection>
<intersection>-118 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-118,36.5,-118</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>474 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-128,41,-128</points>
<connection>
<GID>18</GID>
<name>OUT_11</name></connection>
<connection>
<GID>59</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>478 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-127,41,-127</points>
<connection>
<GID>18</GID>
<name>OUT_12</name></connection>
<connection>
<GID>59</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>470 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-126,41,-126</points>
<connection>
<GID>18</GID>
<name>OUT_13</name></connection>
<connection>
<GID>59</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>472 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-125,41,-125</points>
<connection>
<GID>18</GID>
<name>OUT_14</name></connection>
<connection>
<GID>59</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>476 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-124,41,-124</points>
<connection>
<GID>18</GID>
<name>OUT_15</name></connection>
<connection>
<GID>59</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>96 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-34,-6,-34</points>
<connection>
<GID>6</GID>
<name>IN_3</name></connection>
<connection>
<GID>27</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>463 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-137,41,-137</points>
<connection>
<GID>18</GID>
<name>OUT_2</name></connection>
<connection>
<GID>59</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>464 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-136,41,-136</points>
<connection>
<GID>18</GID>
<name>OUT_3</name></connection>
<connection>
<GID>59</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>466 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-135,41,-135</points>
<connection>
<GID>18</GID>
<name>OUT_4</name></connection>
<connection>
<GID>59</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>468 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-132,41,-132</points>
<connection>
<GID>18</GID>
<name>OUT_7</name></connection>
<connection>
<GID>59</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-7,23,-3</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>-7 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-24.5,-163,-24.5,-7</points>
<intersection>-163 8</intersection>
<intersection>-144 16</intersection>
<intersection>-131.5 34</intersection>
<intersection>-111.5 37</intersection>
<intersection>-70.5 48</intersection>
<intersection>-51 6</intersection>
<intersection>-29.5 55</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24.5,-7,23,-7</points>
<intersection>-24.5 1</intersection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-24.5,-51,22.5,-51</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-24.5,-163,67.5,-163</points>
<intersection>-24.5 1</intersection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-24.5,-144,-13.5,-144</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>67.5,-163,67.5,-29.5</points>
<intersection>-163 8</intersection>
<intersection>-131.5 39</intersection>
<intersection>-111.5 38</intersection>
<intersection>-90 44</intersection>
<intersection>-70.5 50</intersection>
<intersection>-51 49</intersection>
<intersection>-29.5 52</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>-24.5,-131.5,26,-131.5</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-24.5,-111.5,-16,-111.5</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>7.5,-111.5,67.5,-111.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>49.5,-131.5,67.5,-131.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>50,-90,67.5,-90</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-24.5,-70.5,-15.5,-70.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>63.5,-51,67.5,-51</points>
<connection>
<GID>137</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>8,-70.5,67.5,-70.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>36.5,-29.5,67.5,-29.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>67.5 33</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>-24.5,-29.5,-17.5,-29.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>391 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-82.5,46,-82.5</points>
<connection>
<GID>55</GID>
<name>OUT_15</name></connection>
<connection>
<GID>56</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>385 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-90.5,46,-90.5</points>
<connection>
<GID>55</GID>
<name>OUT_7</name></connection>
<connection>
<GID>56</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>389 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-86.5,46,-86.5</points>
<connection>
<GID>55</GID>
<name>OUT_11</name></connection>
<connection>
<GID>56</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>357 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-67,4,-67</points>
<connection>
<GID>53</GID>
<name>OUT_11</name></connection>
<connection>
<GID>54</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>384 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-87.5,46,-87.5</points>
<connection>
<GID>55</GID>
<name>OUT_10</name></connection>
<connection>
<GID>56</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>353 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-71,4,-71</points>
<connection>
<GID>53</GID>
<name>OUT_7</name></connection>
<connection>
<GID>54</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>694 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-61.5,1.5,-59.5</points>
<connection>
<GID>53</GID>
<name>ENABLE_0</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1.5,-59.5,6,-59.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>365 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-78,4,-78</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<connection>
<GID>54</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>366 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-77,4,-77</points>
<connection>
<GID>53</GID>
<name>OUT_1</name></connection>
<connection>
<GID>54</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>351 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-66,4,-66</points>
<connection>
<GID>53</GID>
<name>OUT_12</name></connection>
<connection>
<GID>54</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-13,3.5,14.5</points>
<intersection>-13 1</intersection>
<intersection>14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-13,15.5,-13</points>
<intersection>3.5 0</intersection>
<intersection>15.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,14.5,8.5,14.5</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>3.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15.5,-29.5,15.5,-13</points>
<intersection>-29.5 4</intersection>
<intersection>-29.5 4</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>11,-29.5,18.5,-29.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>15.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>358 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-65,4,-65</points>
<connection>
<GID>53</GID>
<name>OUT_13</name></connection>
<connection>
<GID>54</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>359 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-63,4,-63</points>
<connection>
<GID>53</GID>
<name>OUT_15</name></connection>
<connection>
<GID>54</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>362 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-76,4,-76</points>
<connection>
<GID>53</GID>
<name>OUT_2</name></connection>
<connection>
<GID>54</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>363 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-75,4,-75</points>
<connection>
<GID>53</GID>
<name>OUT_3</name></connection>
<connection>
<GID>54</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>696 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-102.5,1,-100.5</points>
<connection>
<GID>57</GID>
<name>ENABLE_0</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-100.5,5,-100.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>361 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-73,4,-73</points>
<connection>
<GID>53</GID>
<name>OUT_5</name></connection>
<connection>
<GID>54</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>203 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,17,14,17</points>
<connection>
<GID>2</GID>
<name>ADDRESS_10</name></connection>
<connection>
<GID>67</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>364 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-72,4,-72</points>
<connection>
<GID>53</GID>
<name>OUT_6</name></connection>
<connection>
<GID>54</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>201 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,10,14,10</points>
<connection>
<GID>2</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>67</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>354 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-70,4,-70</points>
<connection>
<GID>53</GID>
<name>OUT_8</name></connection>
<connection>
<GID>54</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>355 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-69,4,-69</points>
<connection>
<GID>53</GID>
<name>OUT_9</name></connection>
<connection>
<GID>54</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>695 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-81,43.5,-79</points>
<connection>
<GID>55</GID>
<name>ENABLE_0</name></connection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-79,49.5,-79</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>397 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-97.5,46,-97.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<connection>
<GID>56</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>398 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-96.5,46,-96.5</points>
<connection>
<GID>55</GID>
<name>OUT_1</name></connection>
<connection>
<GID>56</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>383 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-85.5,46,-85.5</points>
<connection>
<GID>55</GID>
<name>OUT_12</name></connection>
<connection>
<GID>56</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>390 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-84.5,46,-84.5</points>
<connection>
<GID>55</GID>
<name>OUT_13</name></connection>
<connection>
<GID>56</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>693 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-46,52.5,-40</points>
<connection>
<GID>100</GID>
<name>ENABLE_0</name></connection>
<intersection>-46 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-40,53.5,-40</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-46,52.5,-46</points>
<intersection>48 8</intersection>
<intersection>52.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>48,-50,48,-46</points>
<connection>
<GID>99</GID>
<name>ENABLE_0</name></connection>
<intersection>-46 2</intersection></vsegment></shape></wire>
<wire>
<ID>388 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-83.5,46,-83.5</points>
<connection>
<GID>55</GID>
<name>OUT_14</name></connection>
<connection>
<GID>56</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>395 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-94.5,46,-94.5</points>
<connection>
<GID>55</GID>
<name>OUT_3</name></connection>
<connection>
<GID>56</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>697 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-122.5,43,-119.5</points>
<connection>
<GID>59</GID>
<name>ENABLE_0</name></connection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>43,-119.5,46,-119.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>392 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-93.5,46,-93.5</points>
<connection>
<GID>55</GID>
<name>OUT_4</name></connection>
<connection>
<GID>56</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>393 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-92.5,46,-92.5</points>
<connection>
<GID>55</GID>
<name>OUT_5</name></connection>
<connection>
<GID>56</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>396 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-91.5,46,-91.5</points>
<connection>
<GID>55</GID>
<name>OUT_6</name></connection>
<connection>
<GID>56</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>387 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-88.5,46,-88.5</points>
<connection>
<GID>55</GID>
<name>OUT_9</name></connection>
<connection>
<GID>56</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>429 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-119,3.5,-119</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<connection>
<GID>58</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>430 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-118,3.5,-118</points>
<connection>
<GID>57</GID>
<name>OUT_1</name></connection>
<connection>
<GID>58</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>416 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-109,3.5,-109</points>
<connection>
<GID>57</GID>
<name>OUT_10</name></connection>
<connection>
<GID>58</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>421 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-108,3.5,-108</points>
<connection>
<GID>57</GID>
<name>OUT_11</name></connection>
<connection>
<GID>58</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>420 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-105,3.5,-105</points>
<connection>
<GID>57</GID>
<name>OUT_14</name></connection>
<connection>
<GID>58</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>426 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-117,3.5,-117</points>
<connection>
<GID>57</GID>
<name>OUT_2</name></connection>
<connection>
<GID>58</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>427 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-116,3.5,-116</points>
<connection>
<GID>57</GID>
<name>OUT_3</name></connection>
<connection>
<GID>58</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>424 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-115,3.5,-115</points>
<connection>
<GID>57</GID>
<name>OUT_4</name></connection>
<connection>
<GID>58</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>425 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-114,3.5,-114</points>
<connection>
<GID>57</GID>
<name>OUT_5</name></connection>
<connection>
<GID>58</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>428 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-113,3.5,-113</points>
<connection>
<GID>57</GID>
<name>OUT_6</name></connection>
<connection>
<GID>58</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>418 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-111,3.5,-111</points>
<connection>
<GID>57</GID>
<name>OUT_8</name></connection>
<connection>
<GID>58</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>419 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-110,3.5,-110</points>
<connection>
<GID>57</GID>
<name>OUT_9</name></connection>
<connection>
<GID>58</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>417 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-112,3.5,-112</points>
<connection>
<GID>57</GID>
<name>OUT_7</name></connection>
<connection>
<GID>58</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>448 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-129,45.5,-129</points>
<connection>
<GID>59</GID>
<name>OUT_10</name></connection>
<connection>
<GID>60</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>94 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-30,-6,-30</points>
<connection>
<GID>6</GID>
<name>IN_7</name></connection>
<connection>
<GID>27</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>453 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-128,45.5,-128</points>
<connection>
<GID>59</GID>
<name>OUT_11</name></connection>
<connection>
<GID>60</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>447 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-127,45.5,-127</points>
<connection>
<GID>59</GID>
<name>OUT_12</name></connection>
<connection>
<GID>60</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>454 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-126,45.5,-126</points>
<connection>
<GID>59</GID>
<name>OUT_13</name></connection>
<connection>
<GID>60</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>452 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-125,45.5,-125</points>
<connection>
<GID>59</GID>
<name>OUT_14</name></connection>
<connection>
<GID>60</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>455 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-124,45.5,-124</points>
<connection>
<GID>59</GID>
<name>OUT_15</name></connection>
<connection>
<GID>60</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>458 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-137,45.5,-137</points>
<connection>
<GID>59</GID>
<name>OUT_2</name></connection>
<connection>
<GID>60</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>456 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-135,45.5,-135</points>
<connection>
<GID>59</GID>
<name>OUT_4</name></connection>
<connection>
<GID>60</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>98 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-32,-6,-32</points>
<connection>
<GID>6</GID>
<name>IN_5</name></connection>
<connection>
<GID>27</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>457 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-134,45.5,-134</points>
<connection>
<GID>59</GID>
<name>OUT_5</name></connection>
<connection>
<GID>60</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>460 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-133,45.5,-133</points>
<connection>
<GID>59</GID>
<name>OUT_6</name></connection>
<connection>
<GID>60</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>449 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-132,45.5,-132</points>
<connection>
<GID>59</GID>
<name>OUT_7</name></connection>
<connection>
<GID>60</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>662 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-57.5,59.5,-57.5</points>
<connection>
<GID>99</GID>
<name>OUT_1</name></connection>
<connection>
<GID>137</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>663 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-56.5,59.5,-56.5</points>
<connection>
<GID>99</GID>
<name>OUT_2</name></connection>
<connection>
<GID>137</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>664 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-55.5,59.5,-55.5</points>
<connection>
<GID>99</GID>
<name>OUT_3</name></connection>
<connection>
<GID>137</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>666 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-53.5,59.5,-53.5</points>
<connection>
<GID>99</GID>
<name>OUT_5</name></connection>
<connection>
<GID>137</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>667 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-52.5,59.5,-52.5</points>
<connection>
<GID>99</GID>
<name>OUT_6</name></connection>
<connection>
<GID>137</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>668 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-51.5,59.5,-51.5</points>
<connection>
<GID>99</GID>
<name>OUT_7</name></connection>
<connection>
<GID>137</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>658 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-49.5,59.5,-49.5</points>
<connection>
<GID>100</GID>
<name>OUT_1</name></connection>
<connection>
<GID>137</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>660 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-48.5,59.5,-48.5</points>
<connection>
<GID>100</GID>
<name>OUT_2</name></connection>
<connection>
<GID>137</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>659 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-47.5,59.5,-47.5</points>
<connection>
<GID>100</GID>
<name>OUT_3</name></connection>
<connection>
<GID>137</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>93 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-35,-6,-35</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<connection>
<GID>27</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>95 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-37,-6,-37</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>97 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-33,-6,-33</points>
<connection>
<GID>6</GID>
<name>IN_4</name></connection>
<connection>
<GID>27</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>175 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-28,-6,-28</points>
<connection>
<GID>6</GID>
<name>IN_9</name></connection>
<connection>
<GID>27</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>176 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-31,-6,-31</points>
<connection>
<GID>6</GID>
<name>IN_6</name></connection>
<connection>
<GID>27</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>177 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-27,-6,-27</points>
<connection>
<GID>6</GID>
<name>IN_10</name></connection>
<connection>
<GID>27</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>178 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-26,-6,-26</points>
<connection>
<GID>6</GID>
<name>IN_11</name></connection>
<connection>
<GID>27</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>179 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-36,-6,-36</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<connection>
<GID>27</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>180 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-29,-6,-29</points>
<connection>
<GID>6</GID>
<name>IN_8</name></connection>
<connection>
<GID>27</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>181 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-33,7,-33</points>
<connection>
<GID>6</GID>
<name>OUT_4</name></connection>
<connection>
<GID>66</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>182 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-36,7,-36</points>
<connection>
<GID>6</GID>
<name>OUT_1</name></connection>
<connection>
<GID>66</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>183 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-32,7,-32</points>
<connection>
<GID>6</GID>
<name>OUT_5</name></connection>
<connection>
<GID>66</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>184 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-31,7,-31</points>
<connection>
<GID>6</GID>
<name>OUT_6</name></connection>
<connection>
<GID>66</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>185 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-30,7,-30</points>
<connection>
<GID>6</GID>
<name>OUT_7</name></connection>
<connection>
<GID>66</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>186 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-28,7,-28</points>
<connection>
<GID>6</GID>
<name>OUT_9</name></connection>
<connection>
<GID>66</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>187 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-29,7,-29</points>
<connection>
<GID>6</GID>
<name>OUT_8</name></connection>
<connection>
<GID>66</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>188 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-37,7,-37</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>189 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-34,7,-34</points>
<connection>
<GID>6</GID>
<name>OUT_3</name></connection>
<connection>
<GID>66</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>190 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-35,7,-35</points>
<connection>
<GID>6</GID>
<name>OUT_2</name></connection>
<connection>
<GID>66</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>191 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-27,7,-27</points>
<connection>
<GID>6</GID>
<name>OUT_10</name></connection>
<connection>
<GID>66</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>192 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-26,7,-26</points>
<connection>
<GID>6</GID>
<name>OUT_11</name></connection>
<connection>
<GID>66</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>193 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,14,14,14</points>
<connection>
<GID>2</GID>
<name>ADDRESS_7</name></connection>
<connection>
<GID>67</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>194 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,15,14,15</points>
<connection>
<GID>2</GID>
<name>ADDRESS_8</name></connection>
<connection>
<GID>67</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>196 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,16,14,16</points>
<connection>
<GID>2</GID>
<name>ADDRESS_9</name></connection>
<connection>
<GID>67</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>197 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,7,14,7</points>
<connection>
<GID>2</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>67</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>198 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,8,14,8</points>
<connection>
<GID>2</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>67</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>199 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,11,14,11</points>
<connection>
<GID>2</GID>
<name>ADDRESS_4</name></connection>
<connection>
<GID>67</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>200 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,13,14,13</points>
<connection>
<GID>2</GID>
<name>ADDRESS_6</name></connection>
<connection>
<GID>67</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>202 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,12,14,12</points>
<connection>
<GID>2</GID>
<name>ADDRESS_5</name></connection>
<connection>
<GID>67</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>204 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,18,14,18</points>
<connection>
<GID>2</GID>
<name>ADDRESS_11</name></connection>
<connection>
<GID>67</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>258 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-93.5,31,-93.5</points>
<connection>
<GID>14</GID>
<name>IN_4</name></connection>
<connection>
<GID>85</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>262 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-85.5,31,-85.5</points>
<connection>
<GID>14</GID>
<name>IN_12</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>266 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-86.5,31,-86.5</points>
<connection>
<GID>14</GID>
<name>IN_11</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>254 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-97.5,31,-97.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>272 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-37,23.5,-37</points>
<connection>
<GID>68</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>255 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-96.5,31,-96.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<connection>
<GID>73</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>257 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-94.5,31,-94.5</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<connection>
<GID>77</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>259 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-91.5,31,-91.5</points>
<connection>
<GID>14</GID>
<name>IN_6</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>261 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-87.5,31,-87.5</points>
<connection>
<GID>14</GID>
<name>IN_10</name></connection>
<connection>
<GID>91</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>263 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-83.5,31,-83.5</points>
<connection>
<GID>14</GID>
<name>IN_14</name></connection>
<connection>
<GID>95</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>265 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-84.5,31,-84.5</points>
<connection>
<GID>14</GID>
<name>IN_13</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>267 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-88.5,31,-88.5</points>
<connection>
<GID>14</GID>
<name>IN_9</name></connection>
<connection>
<GID>90</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>269 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-92.5,31,-92.5</points>
<connection>
<GID>14</GID>
<name>IN_5</name></connection>
<connection>
<GID>86</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>271 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-32,23.5,-32</points>
<connection>
<GID>68</GID>
<name>IN_5</name></connection>
<connection>
<GID>101</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>273 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-35,23.5,-35</points>
<connection>
<GID>68</GID>
<name>IN_2</name></connection>
<connection>
<GID>101</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>274 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-31,23.5,-31</points>
<connection>
<GID>68</GID>
<name>IN_6</name></connection>
<connection>
<GID>101</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>275 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-34,23.5,-34</points>
<connection>
<GID>68</GID>
<name>IN_3</name></connection>
<connection>
<GID>101</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>276 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-36,23.5,-36</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<connection>
<GID>101</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>278 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22.5,-30,23.5,-30</points>
<connection>
<GID>68</GID>
<name>IN_7</name></connection>
<connection>
<GID>101</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>279 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32,-29,32.5,-29</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>280 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32,-28,32.5,-28</points>
<connection>
<GID>102</GID>
<name>OUT_1</name></connection>
<connection>
<GID>24</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>282 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32,-27,32.5,-27</points>
<connection>
<GID>102</GID>
<name>OUT_2</name></connection>
<connection>
<GID>24</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>283 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-29,28,-29</points>
<connection>
<GID>68</GID>
<name>IN_8</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>284 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-28,28,-28</points>
<connection>
<GID>68</GID>
<name>IN_9</name></connection>
<connection>
<GID>102</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>285 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-27,28,-27</points>
<connection>
<GID>68</GID>
<name>IN_10</name></connection>
<connection>
<GID>102</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>286 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-26,28,-26</points>
<connection>
<GID>68</GID>
<name>IN_11</name></connection>
<connection>
<GID>102</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>287 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-30,32.5,-30</points>
<connection>
<GID>101</GID>
<name>OUT_7</name></connection>
<connection>
<GID>24</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>289 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-32,32.5,-32</points>
<connection>
<GID>101</GID>
<name>OUT_5</name></connection>
<connection>
<GID>24</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>290 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-33,32.5,-33</points>
<connection>
<GID>101</GID>
<name>OUT_4</name></connection>
<connection>
<GID>24</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>291 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-34,32.5,-34</points>
<connection>
<GID>101</GID>
<name>OUT_3</name></connection>
<connection>
<GID>24</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>292 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-35,32.5,-35</points>
<connection>
<GID>101</GID>
<name>OUT_2</name></connection>
<connection>
<GID>24</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>293 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-36,32.5,-36</points>
<connection>
<GID>101</GID>
<name>OUT_1</name></connection>
<connection>
<GID>24</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>294 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-37,32.5,-37</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>295 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-24.5,30,-18</points>
<connection>
<GID>102</GID>
<name>ENABLE_0</name></connection>
<intersection>-24.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-18,31,-18</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-24.5,30,-24.5</points>
<intersection>25.5 3</intersection>
<intersection>30 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25.5,-28.5,25.5,-24.5</points>
<connection>
<GID>101</GID>
<name>ENABLE_0</name></connection>
<intersection>-24.5 2</intersection></vsegment></shape></wire></page 0></circuit>